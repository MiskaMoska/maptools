localparam input_mask_0_0 = 5'b00001;
localparam input_mask_1_0 = 5'b00001;
localparam input_mask_2_0 = 5'b00001;
localparam input_mask_0_1 = 5'b01101;
localparam input_mask_1_1 = 5'b11101;
localparam input_mask_2_1 = 5'b01001;
localparam input_mask_0_2 = 5'b01000;
localparam input_mask_1_2 = 5'b00101;
localparam input_mask_2_2 = 5'b00001;

localparam output_sel_0_0 = 5'b10000;
localparam output_sel_1_0 = 5'b10000;
localparam output_sel_2_0 = 5'b10000;
localparam output_sel_0_1 = 5'b10000;
localparam output_sel_1_1 = 5'b00010;
localparam output_sel_2_1 = 5'b00010;
localparam output_sel_0_2 = 5'b00001;
localparam output_sel_1_2 = 5'b01000;
localparam output_sel_2_2 = 5'b00010;