`include "params.svh"
`include "network_config.svh"

module network(
    input       wire                        clk,
    input       wire                        rstn,

    //stab port
    input       wire        [`DW-1:0]       data_i_stab,
    input       wire                        valid_i_stab,
    output      wire                        ready_o_stab,

    //flee0 port
    output      wire        [`DW-1:0]       data_o_flee0,
    output      wire                        valid_o_flee0,
    input       wire                        ready_i_flee0,

    //flee1 port
    output      wire        [`DW-1:0]       data_o_flee1,
    output      wire                        valid_o_flee1,
    input       wire                        ready_i_flee1,

    input       wire        [`DW-1:0]       cast_data_i_0_0,
    input       wire                        cast_valid_i_0_0,
    output      wire                        cast_ready_o_0_0,

    output      wire        [`DW-1:0]       cast_data_o_0_0,
    output      wire                        cast_valid_o_0_0,
    input       wire                        cast_ready_i_0_0,

    input       wire        [`DW-1:0]       cast_data_i_0_1,
    input       wire                        cast_valid_i_0_1,
    output      wire                        cast_ready_o_0_1,

    output      wire        [`DW-1:0]       cast_data_o_0_1,
    output      wire                        cast_valid_o_0_1,
    input       wire                        cast_ready_i_0_1,

    input       wire        [`DW-1:0]       cast_data_i_0_2,
    input       wire                        cast_valid_i_0_2,
    output      wire                        cast_ready_o_0_2,

    output      wire        [`DW-1:0]       cast_data_o_0_2,
    output      wire                        cast_valid_o_0_2,
    input       wire                        cast_ready_i_0_2,

    input       wire        [`DW-1:0]       cast_data_i_0_3,
    input       wire                        cast_valid_i_0_3,
    output      wire                        cast_ready_o_0_3,

    output      wire        [`DW-1:0]       cast_data_o_0_3,
    output      wire                        cast_valid_o_0_3,
    input       wire                        cast_ready_i_0_3,

    input       wire        [`DW-1:0]       cast_data_i_0_4,
    input       wire                        cast_valid_i_0_4,
    output      wire                        cast_ready_o_0_4,

    output      wire        [`DW-1:0]       cast_data_o_0_4,
    output      wire                        cast_valid_o_0_4,
    input       wire                        cast_ready_i_0_4,

    input       wire        [`DW-1:0]       cast_data_i_0_5,
    input       wire                        cast_valid_i_0_5,
    output      wire                        cast_ready_o_0_5,

    output      wire        [`DW-1:0]       cast_data_o_0_5,
    output      wire                        cast_valid_o_0_5,
    input       wire                        cast_ready_i_0_5,

    input       wire        [`DW-1:0]       cast_data_i_0_6,
    input       wire                        cast_valid_i_0_6,
    output      wire                        cast_ready_o_0_6,

    output      wire        [`DW-1:0]       cast_data_o_0_6,
    output      wire                        cast_valid_o_0_6,
    input       wire                        cast_ready_i_0_6,

    input       wire        [`DW-1:0]       cast_data_i_0_7,
    input       wire                        cast_valid_i_0_7,
    output      wire                        cast_ready_o_0_7,

    output      wire        [`DW-1:0]       cast_data_o_0_7,
    output      wire                        cast_valid_o_0_7,
    input       wire                        cast_ready_i_0_7,

    input       wire        [`DW-1:0]       cast_data_i_0_8,
    input       wire                        cast_valid_i_0_8,
    output      wire                        cast_ready_o_0_8,

    output      wire        [`DW-1:0]       cast_data_o_0_8,
    output      wire                        cast_valid_o_0_8,
    input       wire                        cast_ready_i_0_8,

    input       wire        [`DW-1:0]       cast_data_i_0_9,
    input       wire                        cast_valid_i_0_9,
    output      wire                        cast_ready_o_0_9,

    output      wire        [`DW-1:0]       cast_data_o_0_9,
    output      wire                        cast_valid_o_0_9,
    input       wire                        cast_ready_i_0_9,

    input       wire        [`DW-1:0]       cast_data_i_1_0,
    input       wire                        cast_valid_i_1_0,
    output      wire                        cast_ready_o_1_0,

    output      wire        [`DW-1:0]       cast_data_o_1_0,
    output      wire                        cast_valid_o_1_0,
    input       wire                        cast_ready_i_1_0,

    input       wire        [`DW-1:0]       cast_data_i_1_1,
    input       wire                        cast_valid_i_1_1,
    output      wire                        cast_ready_o_1_1,

    output      wire        [`DW-1:0]       cast_data_o_1_1,
    output      wire                        cast_valid_o_1_1,
    input       wire                        cast_ready_i_1_1,

    input       wire        [`DW-1:0]       cast_data_i_1_2,
    input       wire                        cast_valid_i_1_2,
    output      wire                        cast_ready_o_1_2,

    output      wire        [`DW-1:0]       cast_data_o_1_2,
    output      wire                        cast_valid_o_1_2,
    input       wire                        cast_ready_i_1_2,

    input       wire        [`DW-1:0]       cast_data_i_1_3,
    input       wire                        cast_valid_i_1_3,
    output      wire                        cast_ready_o_1_3,

    output      wire        [`DW-1:0]       cast_data_o_1_3,
    output      wire                        cast_valid_o_1_3,
    input       wire                        cast_ready_i_1_3,

    input       wire        [`DW-1:0]       cast_data_i_1_4,
    input       wire                        cast_valid_i_1_4,
    output      wire                        cast_ready_o_1_4,

    output      wire        [`DW-1:0]       cast_data_o_1_4,
    output      wire                        cast_valid_o_1_4,
    input       wire                        cast_ready_i_1_4,

    input       wire        [`DW-1:0]       cast_data_i_1_5,
    input       wire                        cast_valid_i_1_5,
    output      wire                        cast_ready_o_1_5,

    output      wire        [`DW-1:0]       cast_data_o_1_5,
    output      wire                        cast_valid_o_1_5,
    input       wire                        cast_ready_i_1_5,

    input       wire        [`DW-1:0]       cast_data_i_1_6,
    input       wire                        cast_valid_i_1_6,
    output      wire                        cast_ready_o_1_6,

    output      wire        [`DW-1:0]       cast_data_o_1_6,
    output      wire                        cast_valid_o_1_6,
    input       wire                        cast_ready_i_1_6,

    input       wire        [`DW-1:0]       cast_data_i_1_7,
    input       wire                        cast_valid_i_1_7,
    output      wire                        cast_ready_o_1_7,

    output      wire        [`DW-1:0]       cast_data_o_1_7,
    output      wire                        cast_valid_o_1_7,
    input       wire                        cast_ready_i_1_7,

    input       wire        [`DW-1:0]       cast_data_i_1_8,
    input       wire                        cast_valid_i_1_8,
    output      wire                        cast_ready_o_1_8,

    output      wire        [`DW-1:0]       cast_data_o_1_8,
    output      wire                        cast_valid_o_1_8,
    input       wire                        cast_ready_i_1_8,

    input       wire        [`DW-1:0]       cast_data_i_1_9,
    input       wire                        cast_valid_i_1_9,
    output      wire                        cast_ready_o_1_9,

    output      wire        [`DW-1:0]       cast_data_o_1_9,
    output      wire                        cast_valid_o_1_9,
    input       wire                        cast_ready_i_1_9,

    input       wire        [`DW-1:0]       cast_data_i_2_0,
    input       wire                        cast_valid_i_2_0,
    output      wire                        cast_ready_o_2_0,

    output      wire        [`DW-1:0]       cast_data_o_2_0,
    output      wire                        cast_valid_o_2_0,
    input       wire                        cast_ready_i_2_0,

    input       wire        [`DW-1:0]       cast_data_i_2_1,
    input       wire                        cast_valid_i_2_1,
    output      wire                        cast_ready_o_2_1,

    output      wire        [`DW-1:0]       cast_data_o_2_1,
    output      wire                        cast_valid_o_2_1,
    input       wire                        cast_ready_i_2_1,

    input       wire        [`DW-1:0]       cast_data_i_2_2,
    input       wire                        cast_valid_i_2_2,
    output      wire                        cast_ready_o_2_2,

    output      wire        [`DW-1:0]       cast_data_o_2_2,
    output      wire                        cast_valid_o_2_2,
    input       wire                        cast_ready_i_2_2,

    input       wire        [`DW-1:0]       cast_data_i_2_3,
    input       wire                        cast_valid_i_2_3,
    output      wire                        cast_ready_o_2_3,

    output      wire        [`DW-1:0]       cast_data_o_2_3,
    output      wire                        cast_valid_o_2_3,
    input       wire                        cast_ready_i_2_3,

    input       wire        [`DW-1:0]       cast_data_i_2_4,
    input       wire                        cast_valid_i_2_4,
    output      wire                        cast_ready_o_2_4,

    output      wire        [`DW-1:0]       cast_data_o_2_4,
    output      wire                        cast_valid_o_2_4,
    input       wire                        cast_ready_i_2_4,

    input       wire        [`DW-1:0]       cast_data_i_2_5,
    input       wire                        cast_valid_i_2_5,
    output      wire                        cast_ready_o_2_5,

    output      wire        [`DW-1:0]       cast_data_o_2_5,
    output      wire                        cast_valid_o_2_5,
    input       wire                        cast_ready_i_2_5,

    input       wire        [`DW-1:0]       cast_data_i_2_6,
    input       wire                        cast_valid_i_2_6,
    output      wire                        cast_ready_o_2_6,

    output      wire        [`DW-1:0]       cast_data_o_2_6,
    output      wire                        cast_valid_o_2_6,
    input       wire                        cast_ready_i_2_6,

    input       wire        [`DW-1:0]       cast_data_i_2_7,
    input       wire                        cast_valid_i_2_7,
    output      wire                        cast_ready_o_2_7,

    output      wire        [`DW-1:0]       cast_data_o_2_7,
    output      wire                        cast_valid_o_2_7,
    input       wire                        cast_ready_i_2_7,

    input       wire        [`DW-1:0]       cast_data_i_2_8,
    input       wire                        cast_valid_i_2_8,
    output      wire                        cast_ready_o_2_8,

    output      wire        [`DW-1:0]       cast_data_o_2_8,
    output      wire                        cast_valid_o_2_8,
    input       wire                        cast_ready_i_2_8,

    input       wire        [`DW-1:0]       cast_data_i_2_9,
    input       wire                        cast_valid_i_2_9,
    output      wire                        cast_ready_o_2_9,

    output      wire        [`DW-1:0]       cast_data_o_2_9,
    output      wire                        cast_valid_o_2_9,
    input       wire                        cast_ready_i_2_9,

    input       wire        [`DW-1:0]       cast_data_i_3_0,
    input       wire                        cast_valid_i_3_0,
    output      wire                        cast_ready_o_3_0,

    output      wire        [`DW-1:0]       cast_data_o_3_0,
    output      wire                        cast_valid_o_3_0,
    input       wire                        cast_ready_i_3_0,

    input       wire        [`DW-1:0]       cast_data_i_3_1,
    input       wire                        cast_valid_i_3_1,
    output      wire                        cast_ready_o_3_1,

    output      wire        [`DW-1:0]       cast_data_o_3_1,
    output      wire                        cast_valid_o_3_1,
    input       wire                        cast_ready_i_3_1,

    input       wire        [`DW-1:0]       cast_data_i_3_2,
    input       wire                        cast_valid_i_3_2,
    output      wire                        cast_ready_o_3_2,

    output      wire        [`DW-1:0]       cast_data_o_3_2,
    output      wire                        cast_valid_o_3_2,
    input       wire                        cast_ready_i_3_2,

    input       wire        [`DW-1:0]       cast_data_i_3_3,
    input       wire                        cast_valid_i_3_3,
    output      wire                        cast_ready_o_3_3,

    output      wire        [`DW-1:0]       cast_data_o_3_3,
    output      wire                        cast_valid_o_3_3,
    input       wire                        cast_ready_i_3_3,

    input       wire        [`DW-1:0]       cast_data_i_3_4,
    input       wire                        cast_valid_i_3_4,
    output      wire                        cast_ready_o_3_4,

    output      wire        [`DW-1:0]       cast_data_o_3_4,
    output      wire                        cast_valid_o_3_4,
    input       wire                        cast_ready_i_3_4,

    input       wire        [`DW-1:0]       cast_data_i_3_5,
    input       wire                        cast_valid_i_3_5,
    output      wire                        cast_ready_o_3_5,

    output      wire        [`DW-1:0]       cast_data_o_3_5,
    output      wire                        cast_valid_o_3_5,
    input       wire                        cast_ready_i_3_5,

    input       wire        [`DW-1:0]       cast_data_i_3_6,
    input       wire                        cast_valid_i_3_6,
    output      wire                        cast_ready_o_3_6,

    output      wire        [`DW-1:0]       cast_data_o_3_6,
    output      wire                        cast_valid_o_3_6,
    input       wire                        cast_ready_i_3_6,

    input       wire        [`DW-1:0]       cast_data_i_3_7,
    input       wire                        cast_valid_i_3_7,
    output      wire                        cast_ready_o_3_7,

    output      wire        [`DW-1:0]       cast_data_o_3_7,
    output      wire                        cast_valid_o_3_7,
    input       wire                        cast_ready_i_3_7,

    input       wire        [`DW-1:0]       cast_data_i_3_8,
    input       wire                        cast_valid_i_3_8,
    output      wire                        cast_ready_o_3_8,

    output      wire        [`DW-1:0]       cast_data_o_3_8,
    output      wire                        cast_valid_o_3_8,
    input       wire                        cast_ready_i_3_8,

    input       wire        [`DW-1:0]       cast_data_i_3_9,
    input       wire                        cast_valid_i_3_9,
    output      wire                        cast_ready_o_3_9,

    output      wire        [`DW-1:0]       cast_data_o_3_9,
    output      wire                        cast_valid_o_3_9,
    input       wire                        cast_ready_i_3_9,

    input       wire        [`DW-1:0]       cast_data_i_4_0,
    input       wire                        cast_valid_i_4_0,
    output      wire                        cast_ready_o_4_0,

    output      wire        [`DW-1:0]       cast_data_o_4_0,
    output      wire                        cast_valid_o_4_0,
    input       wire                        cast_ready_i_4_0,

    input       wire        [`DW-1:0]       cast_data_i_4_1,
    input       wire                        cast_valid_i_4_1,
    output      wire                        cast_ready_o_4_1,

    output      wire        [`DW-1:0]       cast_data_o_4_1,
    output      wire                        cast_valid_o_4_1,
    input       wire                        cast_ready_i_4_1,

    input       wire        [`DW-1:0]       cast_data_i_4_2,
    input       wire                        cast_valid_i_4_2,
    output      wire                        cast_ready_o_4_2,

    output      wire        [`DW-1:0]       cast_data_o_4_2,
    output      wire                        cast_valid_o_4_2,
    input       wire                        cast_ready_i_4_2,

    input       wire        [`DW-1:0]       cast_data_i_4_3,
    input       wire                        cast_valid_i_4_3,
    output      wire                        cast_ready_o_4_3,

    output      wire        [`DW-1:0]       cast_data_o_4_3,
    output      wire                        cast_valid_o_4_3,
    input       wire                        cast_ready_i_4_3,

    input       wire        [`DW-1:0]       cast_data_i_4_4,
    input       wire                        cast_valid_i_4_4,
    output      wire                        cast_ready_o_4_4,

    output      wire        [`DW-1:0]       cast_data_o_4_4,
    output      wire                        cast_valid_o_4_4,
    input       wire                        cast_ready_i_4_4,

    input       wire        [`DW-1:0]       cast_data_i_4_5,
    input       wire                        cast_valid_i_4_5,
    output      wire                        cast_ready_o_4_5,

    output      wire        [`DW-1:0]       cast_data_o_4_5,
    output      wire                        cast_valid_o_4_5,
    input       wire                        cast_ready_i_4_5,

    input       wire        [`DW-1:0]       cast_data_i_4_6,
    input       wire                        cast_valid_i_4_6,
    output      wire                        cast_ready_o_4_6,

    output      wire        [`DW-1:0]       cast_data_o_4_6,
    output      wire                        cast_valid_o_4_6,
    input       wire                        cast_ready_i_4_6,

    input       wire        [`DW-1:0]       cast_data_i_4_7,
    input       wire                        cast_valid_i_4_7,
    output      wire                        cast_ready_o_4_7,

    output      wire        [`DW-1:0]       cast_data_o_4_7,
    output      wire                        cast_valid_o_4_7,
    input       wire                        cast_ready_i_4_7,

    input       wire        [`DW-1:0]       cast_data_i_4_8,
    input       wire                        cast_valid_i_4_8,
    output      wire                        cast_ready_o_4_8,

    output      wire        [`DW-1:0]       cast_data_o_4_8,
    output      wire                        cast_valid_o_4_8,
    input       wire                        cast_ready_i_4_8,

    input       wire        [`DW-1:0]       cast_data_i_4_9,
    input       wire                        cast_valid_i_4_9,
    output      wire                        cast_ready_o_4_9,

    output      wire        [`DW-1:0]       cast_data_o_4_9,
    output      wire                        cast_valid_o_4_9,
    input       wire                        cast_ready_i_4_9,

    input       wire        [`DW-1:0]       merge_data_i_0_0,
    input       wire                        merge_valid_i_0_0,
    output      wire                        merge_ready_o_0_0,

    output      wire        [`DW-1:0]       merge_data_o_0_0,
    output      wire                        merge_valid_o_0_0,
    input       wire                        merge_ready_i_0_0,
    input       wire        [`DW-1:0]       merge_data_i_0_1,
    input       wire                        merge_valid_i_0_1,
    output      wire                        merge_ready_o_0_1,

    output      wire        [`DW-1:0]       merge_data_o_0_1,
    output      wire                        merge_valid_o_0_1,
    input       wire                        merge_ready_i_0_1,
    input       wire        [`DW-1:0]       merge_data_i_0_2,
    input       wire                        merge_valid_i_0_2,
    output      wire                        merge_ready_o_0_2,

    output      wire        [`DW-1:0]       merge_data_o_0_2,
    output      wire                        merge_valid_o_0_2,
    input       wire                        merge_ready_i_0_2,
    input       wire        [`DW-1:0]       merge_data_i_0_3,
    input       wire                        merge_valid_i_0_3,
    output      wire                        merge_ready_o_0_3,

    output      wire        [`DW-1:0]       merge_data_o_0_3,
    output      wire                        merge_valid_o_0_3,
    input       wire                        merge_ready_i_0_3,
    input       wire        [`DW-1:0]       merge_data_i_0_4,
    input       wire                        merge_valid_i_0_4,
    output      wire                        merge_ready_o_0_4,

    output      wire        [`DW-1:0]       merge_data_o_0_4,
    output      wire                        merge_valid_o_0_4,
    input       wire                        merge_ready_i_0_4,
    input       wire        [`DW-1:0]       merge_data_i_0_5,
    input       wire                        merge_valid_i_0_5,
    output      wire                        merge_ready_o_0_5,

    output      wire        [`DW-1:0]       merge_data_o_0_5,
    output      wire                        merge_valid_o_0_5,
    input       wire                        merge_ready_i_0_5,
    input       wire        [`DW-1:0]       merge_data_i_0_6,
    input       wire                        merge_valid_i_0_6,
    output      wire                        merge_ready_o_0_6,

    output      wire        [`DW-1:0]       merge_data_o_0_6,
    output      wire                        merge_valid_o_0_6,
    input       wire                        merge_ready_i_0_6,
    input       wire        [`DW-1:0]       merge_data_i_0_7,
    input       wire                        merge_valid_i_0_7,
    output      wire                        merge_ready_o_0_7,

    output      wire        [`DW-1:0]       merge_data_o_0_7,
    output      wire                        merge_valid_o_0_7,
    input       wire                        merge_ready_i_0_7,
    input       wire        [`DW-1:0]       merge_data_i_0_8,
    input       wire                        merge_valid_i_0_8,
    output      wire                        merge_ready_o_0_8,

    output      wire        [`DW-1:0]       merge_data_o_0_8,
    output      wire                        merge_valid_o_0_8,
    input       wire                        merge_ready_i_0_8,
    input       wire        [`DW-1:0]       merge_data_i_0_9,
    input       wire                        merge_valid_i_0_9,
    output      wire                        merge_ready_o_0_9,

    output      wire        [`DW-1:0]       merge_data_o_0_9,
    output      wire                        merge_valid_o_0_9,
    input       wire                        merge_ready_i_0_9,
    input       wire        [`DW-1:0]       merge_data_i_1_0,
    input       wire                        merge_valid_i_1_0,
    output      wire                        merge_ready_o_1_0,

    output      wire        [`DW-1:0]       merge_data_o_1_0,
    output      wire                        merge_valid_o_1_0,
    input       wire                        merge_ready_i_1_0,
    input       wire        [`DW-1:0]       merge_data_i_1_1,
    input       wire                        merge_valid_i_1_1,
    output      wire                        merge_ready_o_1_1,

    output      wire        [`DW-1:0]       merge_data_o_1_1,
    output      wire                        merge_valid_o_1_1,
    input       wire                        merge_ready_i_1_1,
    input       wire        [`DW-1:0]       merge_data_i_1_2,
    input       wire                        merge_valid_i_1_2,
    output      wire                        merge_ready_o_1_2,

    output      wire        [`DW-1:0]       merge_data_o_1_2,
    output      wire                        merge_valid_o_1_2,
    input       wire                        merge_ready_i_1_2,
    input       wire        [`DW-1:0]       merge_data_i_1_3,
    input       wire                        merge_valid_i_1_3,
    output      wire                        merge_ready_o_1_3,

    output      wire        [`DW-1:0]       merge_data_o_1_3,
    output      wire                        merge_valid_o_1_3,
    input       wire                        merge_ready_i_1_3,
    input       wire        [`DW-1:0]       merge_data_i_1_4,
    input       wire                        merge_valid_i_1_4,
    output      wire                        merge_ready_o_1_4,

    output      wire        [`DW-1:0]       merge_data_o_1_4,
    output      wire                        merge_valid_o_1_4,
    input       wire                        merge_ready_i_1_4,
    input       wire        [`DW-1:0]       merge_data_i_1_5,
    input       wire                        merge_valid_i_1_5,
    output      wire                        merge_ready_o_1_5,

    output      wire        [`DW-1:0]       merge_data_o_1_5,
    output      wire                        merge_valid_o_1_5,
    input       wire                        merge_ready_i_1_5,
    input       wire        [`DW-1:0]       merge_data_i_1_6,
    input       wire                        merge_valid_i_1_6,
    output      wire                        merge_ready_o_1_6,

    output      wire        [`DW-1:0]       merge_data_o_1_6,
    output      wire                        merge_valid_o_1_6,
    input       wire                        merge_ready_i_1_6,
    input       wire        [`DW-1:0]       merge_data_i_1_7,
    input       wire                        merge_valid_i_1_7,
    output      wire                        merge_ready_o_1_7,

    output      wire        [`DW-1:0]       merge_data_o_1_7,
    output      wire                        merge_valid_o_1_7,
    input       wire                        merge_ready_i_1_7,
    input       wire        [`DW-1:0]       merge_data_i_1_8,
    input       wire                        merge_valid_i_1_8,
    output      wire                        merge_ready_o_1_8,

    output      wire        [`DW-1:0]       merge_data_o_1_8,
    output      wire                        merge_valid_o_1_8,
    input       wire                        merge_ready_i_1_8,
    input       wire        [`DW-1:0]       merge_data_i_1_9,
    input       wire                        merge_valid_i_1_9,
    output      wire                        merge_ready_o_1_9,

    output      wire        [`DW-1:0]       merge_data_o_1_9,
    output      wire                        merge_valid_o_1_9,
    input       wire                        merge_ready_i_1_9,
    input       wire        [`DW-1:0]       merge_data_i_2_0,
    input       wire                        merge_valid_i_2_0,
    output      wire                        merge_ready_o_2_0,

    output      wire        [`DW-1:0]       merge_data_o_2_0,
    output      wire                        merge_valid_o_2_0,
    input       wire                        merge_ready_i_2_0,
    input       wire        [`DW-1:0]       merge_data_i_2_1,
    input       wire                        merge_valid_i_2_1,
    output      wire                        merge_ready_o_2_1,

    output      wire        [`DW-1:0]       merge_data_o_2_1,
    output      wire                        merge_valid_o_2_1,
    input       wire                        merge_ready_i_2_1,
    input       wire        [`DW-1:0]       merge_data_i_2_2,
    input       wire                        merge_valid_i_2_2,
    output      wire                        merge_ready_o_2_2,

    output      wire        [`DW-1:0]       merge_data_o_2_2,
    output      wire                        merge_valid_o_2_2,
    input       wire                        merge_ready_i_2_2,
    input       wire        [`DW-1:0]       merge_data_i_2_3,
    input       wire                        merge_valid_i_2_3,
    output      wire                        merge_ready_o_2_3,

    output      wire        [`DW-1:0]       merge_data_o_2_3,
    output      wire                        merge_valid_o_2_3,
    input       wire                        merge_ready_i_2_3,
    input       wire        [`DW-1:0]       merge_data_i_2_4,
    input       wire                        merge_valid_i_2_4,
    output      wire                        merge_ready_o_2_4,

    output      wire        [`DW-1:0]       merge_data_o_2_4,
    output      wire                        merge_valid_o_2_4,
    input       wire                        merge_ready_i_2_4,
    input       wire        [`DW-1:0]       merge_data_i_2_5,
    input       wire                        merge_valid_i_2_5,
    output      wire                        merge_ready_o_2_5,

    output      wire        [`DW-1:0]       merge_data_o_2_5,
    output      wire                        merge_valid_o_2_5,
    input       wire                        merge_ready_i_2_5,
    input       wire        [`DW-1:0]       merge_data_i_2_6,
    input       wire                        merge_valid_i_2_6,
    output      wire                        merge_ready_o_2_6,

    output      wire        [`DW-1:0]       merge_data_o_2_6,
    output      wire                        merge_valid_o_2_6,
    input       wire                        merge_ready_i_2_6,
    input       wire        [`DW-1:0]       merge_data_i_2_7,
    input       wire                        merge_valid_i_2_7,
    output      wire                        merge_ready_o_2_7,

    output      wire        [`DW-1:0]       merge_data_o_2_7,
    output      wire                        merge_valid_o_2_7,
    input       wire                        merge_ready_i_2_7,
    input       wire        [`DW-1:0]       merge_data_i_2_8,
    input       wire                        merge_valid_i_2_8,
    output      wire                        merge_ready_o_2_8,

    output      wire        [`DW-1:0]       merge_data_o_2_8,
    output      wire                        merge_valid_o_2_8,
    input       wire                        merge_ready_i_2_8,
    input       wire        [`DW-1:0]       merge_data_i_2_9,
    input       wire                        merge_valid_i_2_9,
    output      wire                        merge_ready_o_2_9,

    output      wire        [`DW-1:0]       merge_data_o_2_9,
    output      wire                        merge_valid_o_2_9,
    input       wire                        merge_ready_i_2_9,
    input       wire        [`DW-1:0]       merge_data_i_3_0,
    input       wire                        merge_valid_i_3_0,
    output      wire                        merge_ready_o_3_0,

    output      wire        [`DW-1:0]       merge_data_o_3_0,
    output      wire                        merge_valid_o_3_0,
    input       wire                        merge_ready_i_3_0,
    input       wire        [`DW-1:0]       merge_data_i_3_1,
    input       wire                        merge_valid_i_3_1,
    output      wire                        merge_ready_o_3_1,

    output      wire        [`DW-1:0]       merge_data_o_3_1,
    output      wire                        merge_valid_o_3_1,
    input       wire                        merge_ready_i_3_1,
    input       wire        [`DW-1:0]       merge_data_i_3_2,
    input       wire                        merge_valid_i_3_2,
    output      wire                        merge_ready_o_3_2,

    output      wire        [`DW-1:0]       merge_data_o_3_2,
    output      wire                        merge_valid_o_3_2,
    input       wire                        merge_ready_i_3_2,
    input       wire        [`DW-1:0]       merge_data_i_3_3,
    input       wire                        merge_valid_i_3_3,
    output      wire                        merge_ready_o_3_3,

    output      wire        [`DW-1:0]       merge_data_o_3_3,
    output      wire                        merge_valid_o_3_3,
    input       wire                        merge_ready_i_3_3,
    input       wire        [`DW-1:0]       merge_data_i_3_4,
    input       wire                        merge_valid_i_3_4,
    output      wire                        merge_ready_o_3_4,

    output      wire        [`DW-1:0]       merge_data_o_3_4,
    output      wire                        merge_valid_o_3_4,
    input       wire                        merge_ready_i_3_4,
    input       wire        [`DW-1:0]       merge_data_i_3_5,
    input       wire                        merge_valid_i_3_5,
    output      wire                        merge_ready_o_3_5,

    output      wire        [`DW-1:0]       merge_data_o_3_5,
    output      wire                        merge_valid_o_3_5,
    input       wire                        merge_ready_i_3_5,
    input       wire        [`DW-1:0]       merge_data_i_3_6,
    input       wire                        merge_valid_i_3_6,
    output      wire                        merge_ready_o_3_6,

    output      wire        [`DW-1:0]       merge_data_o_3_6,
    output      wire                        merge_valid_o_3_6,
    input       wire                        merge_ready_i_3_6,
    input       wire        [`DW-1:0]       merge_data_i_3_7,
    input       wire                        merge_valid_i_3_7,
    output      wire                        merge_ready_o_3_7,

    output      wire        [`DW-1:0]       merge_data_o_3_7,
    output      wire                        merge_valid_o_3_7,
    input       wire                        merge_ready_i_3_7,
    input       wire        [`DW-1:0]       merge_data_i_3_8,
    input       wire                        merge_valid_i_3_8,
    output      wire                        merge_ready_o_3_8,

    output      wire        [`DW-1:0]       merge_data_o_3_8,
    output      wire                        merge_valid_o_3_8,
    input       wire                        merge_ready_i_3_8,
    input       wire        [`DW-1:0]       merge_data_i_3_9,
    input       wire                        merge_valid_i_3_9,
    output      wire                        merge_ready_o_3_9,

    output      wire        [`DW-1:0]       merge_data_o_3_9,
    output      wire                        merge_valid_o_3_9,
    input       wire                        merge_ready_i_3_9,
    input       wire        [`DW-1:0]       merge_data_i_4_0,
    input       wire                        merge_valid_i_4_0,
    output      wire                        merge_ready_o_4_0,

    output      wire        [`DW-1:0]       merge_data_o_4_0,
    output      wire                        merge_valid_o_4_0,
    input       wire                        merge_ready_i_4_0,
    input       wire        [`DW-1:0]       merge_data_i_4_1,
    input       wire                        merge_valid_i_4_1,
    output      wire                        merge_ready_o_4_1,

    output      wire        [`DW-1:0]       merge_data_o_4_1,
    output      wire                        merge_valid_o_4_1,
    input       wire                        merge_ready_i_4_1,
    input       wire        [`DW-1:0]       merge_data_i_4_2,
    input       wire                        merge_valid_i_4_2,
    output      wire                        merge_ready_o_4_2,

    output      wire        [`DW-1:0]       merge_data_o_4_2,
    output      wire                        merge_valid_o_4_2,
    input       wire                        merge_ready_i_4_2,
    input       wire        [`DW-1:0]       merge_data_i_4_3,
    input       wire                        merge_valid_i_4_3,
    output      wire                        merge_ready_o_4_3,

    output      wire        [`DW-1:0]       merge_data_o_4_3,
    output      wire                        merge_valid_o_4_3,
    input       wire                        merge_ready_i_4_3,
    input       wire        [`DW-1:0]       merge_data_i_4_4,
    input       wire                        merge_valid_i_4_4,
    output      wire                        merge_ready_o_4_4,

    output      wire        [`DW-1:0]       merge_data_o_4_4,
    output      wire                        merge_valid_o_4_4,
    input       wire                        merge_ready_i_4_4,
    input       wire        [`DW-1:0]       merge_data_i_4_5,
    input       wire                        merge_valid_i_4_5,
    output      wire                        merge_ready_o_4_5,

    output      wire        [`DW-1:0]       merge_data_o_4_5,
    output      wire                        merge_valid_o_4_5,
    input       wire                        merge_ready_i_4_5,
    input       wire        [`DW-1:0]       merge_data_i_4_6,
    input       wire                        merge_valid_i_4_6,
    output      wire                        merge_ready_o_4_6,

    output      wire        [`DW-1:0]       merge_data_o_4_6,
    output      wire                        merge_valid_o_4_6,
    input       wire                        merge_ready_i_4_6,
    input       wire        [`DW-1:0]       merge_data_i_4_7,
    input       wire                        merge_valid_i_4_7,
    output      wire                        merge_ready_o_4_7,

    output      wire        [`DW-1:0]       merge_data_o_4_7,
    output      wire                        merge_valid_o_4_7,
    input       wire                        merge_ready_i_4_7,
    input       wire        [`DW-1:0]       merge_data_i_4_8,
    input       wire                        merge_valid_i_4_8,
    output      wire                        merge_ready_o_4_8,

    output      wire        [`DW-1:0]       merge_data_o_4_8,
    output      wire                        merge_valid_o_4_8,
    input       wire                        merge_ready_i_4_8,
    input       wire        [`DW-1:0]       merge_data_i_4_9,
    input       wire                        merge_valid_i_4_9,
    output      wire                        merge_ready_o_4_9,

    output      wire        [`DW-1:0]       merge_data_o_4_9,
    output      wire                        merge_valid_o_4_9,
    input       wire                        merge_ready_i_4_9,
    input       wire        [`DW-1:0]       gather_data_i_0_0,
    input       wire                        gather_valid_i_0_0,
    output      wire                        gather_ready_o_0_0,

    output      wire        [`DW-1:0]       gather_data_o_0_0,
    output      wire                        gather_valid_o_0_0,
    input       wire                        gather_ready_i_0_0,
    input       wire        [`DW-1:0]       gather_data_i_0_1,
    input       wire                        gather_valid_i_0_1,
    output      wire                        gather_ready_o_0_1,

    output      wire        [`DW-1:0]       gather_data_o_0_1,
    output      wire                        gather_valid_o_0_1,
    input       wire                        gather_ready_i_0_1,
    input       wire        [`DW-1:0]       gather_data_i_0_2,
    input       wire                        gather_valid_i_0_2,
    output      wire                        gather_ready_o_0_2,

    output      wire        [`DW-1:0]       gather_data_o_0_2,
    output      wire                        gather_valid_o_0_2,
    input       wire                        gather_ready_i_0_2,
    input       wire        [`DW-1:0]       gather_data_i_0_3,
    input       wire                        gather_valid_i_0_3,
    output      wire                        gather_ready_o_0_3,

    output      wire        [`DW-1:0]       gather_data_o_0_3,
    output      wire                        gather_valid_o_0_3,
    input       wire                        gather_ready_i_0_3,
    input       wire        [`DW-1:0]       gather_data_i_0_4,
    input       wire                        gather_valid_i_0_4,
    output      wire                        gather_ready_o_0_4,

    output      wire        [`DW-1:0]       gather_data_o_0_4,
    output      wire                        gather_valid_o_0_4,
    input       wire                        gather_ready_i_0_4,
    input       wire        [`DW-1:0]       gather_data_i_0_5,
    input       wire                        gather_valid_i_0_5,
    output      wire                        gather_ready_o_0_5,

    output      wire        [`DW-1:0]       gather_data_o_0_5,
    output      wire                        gather_valid_o_0_5,
    input       wire                        gather_ready_i_0_5,
    input       wire        [`DW-1:0]       gather_data_i_0_6,
    input       wire                        gather_valid_i_0_6,
    output      wire                        gather_ready_o_0_6,

    output      wire        [`DW-1:0]       gather_data_o_0_6,
    output      wire                        gather_valid_o_0_6,
    input       wire                        gather_ready_i_0_6,
    input       wire        [`DW-1:0]       gather_data_i_0_7,
    input       wire                        gather_valid_i_0_7,
    output      wire                        gather_ready_o_0_7,

    output      wire        [`DW-1:0]       gather_data_o_0_7,
    output      wire                        gather_valid_o_0_7,
    input       wire                        gather_ready_i_0_7,
    input       wire        [`DW-1:0]       gather_data_i_0_8,
    input       wire                        gather_valid_i_0_8,
    output      wire                        gather_ready_o_0_8,

    output      wire        [`DW-1:0]       gather_data_o_0_8,
    output      wire                        gather_valid_o_0_8,
    input       wire                        gather_ready_i_0_8,
    input       wire        [`DW-1:0]       gather_data_i_0_9,
    input       wire                        gather_valid_i_0_9,
    output      wire                        gather_ready_o_0_9,

    output      wire        [`DW-1:0]       gather_data_o_0_9,
    output      wire                        gather_valid_o_0_9,
    input       wire                        gather_ready_i_0_9,
    input       wire        [`DW-1:0]       gather_data_i_1_0,
    input       wire                        gather_valid_i_1_0,
    output      wire                        gather_ready_o_1_0,

    output      wire        [`DW-1:0]       gather_data_o_1_0,
    output      wire                        gather_valid_o_1_0,
    input       wire                        gather_ready_i_1_0,
    input       wire        [`DW-1:0]       gather_data_i_1_1,
    input       wire                        gather_valid_i_1_1,
    output      wire                        gather_ready_o_1_1,

    output      wire        [`DW-1:0]       gather_data_o_1_1,
    output      wire                        gather_valid_o_1_1,
    input       wire                        gather_ready_i_1_1,
    input       wire        [`DW-1:0]       gather_data_i_1_2,
    input       wire                        gather_valid_i_1_2,
    output      wire                        gather_ready_o_1_2,

    output      wire        [`DW-1:0]       gather_data_o_1_2,
    output      wire                        gather_valid_o_1_2,
    input       wire                        gather_ready_i_1_2,
    input       wire        [`DW-1:0]       gather_data_i_1_3,
    input       wire                        gather_valid_i_1_3,
    output      wire                        gather_ready_o_1_3,

    output      wire        [`DW-1:0]       gather_data_o_1_3,
    output      wire                        gather_valid_o_1_3,
    input       wire                        gather_ready_i_1_3,
    input       wire        [`DW-1:0]       gather_data_i_1_4,
    input       wire                        gather_valid_i_1_4,
    output      wire                        gather_ready_o_1_4,

    output      wire        [`DW-1:0]       gather_data_o_1_4,
    output      wire                        gather_valid_o_1_4,
    input       wire                        gather_ready_i_1_4,
    input       wire        [`DW-1:0]       gather_data_i_1_5,
    input       wire                        gather_valid_i_1_5,
    output      wire                        gather_ready_o_1_5,

    output      wire        [`DW-1:0]       gather_data_o_1_5,
    output      wire                        gather_valid_o_1_5,
    input       wire                        gather_ready_i_1_5,
    input       wire        [`DW-1:0]       gather_data_i_1_6,
    input       wire                        gather_valid_i_1_6,
    output      wire                        gather_ready_o_1_6,

    output      wire        [`DW-1:0]       gather_data_o_1_6,
    output      wire                        gather_valid_o_1_6,
    input       wire                        gather_ready_i_1_6,
    input       wire        [`DW-1:0]       gather_data_i_1_7,
    input       wire                        gather_valid_i_1_7,
    output      wire                        gather_ready_o_1_7,

    output      wire        [`DW-1:0]       gather_data_o_1_7,
    output      wire                        gather_valid_o_1_7,
    input       wire                        gather_ready_i_1_7,
    input       wire        [`DW-1:0]       gather_data_i_1_8,
    input       wire                        gather_valid_i_1_8,
    output      wire                        gather_ready_o_1_8,

    output      wire        [`DW-1:0]       gather_data_o_1_8,
    output      wire                        gather_valid_o_1_8,
    input       wire                        gather_ready_i_1_8,
    input       wire        [`DW-1:0]       gather_data_i_1_9,
    input       wire                        gather_valid_i_1_9,
    output      wire                        gather_ready_o_1_9,

    output      wire        [`DW-1:0]       gather_data_o_1_9,
    output      wire                        gather_valid_o_1_9,
    input       wire                        gather_ready_i_1_9,
    input       wire        [`DW-1:0]       gather_data_i_2_0,
    input       wire                        gather_valid_i_2_0,
    output      wire                        gather_ready_o_2_0,

    output      wire        [`DW-1:0]       gather_data_o_2_0,
    output      wire                        gather_valid_o_2_0,
    input       wire                        gather_ready_i_2_0,
    input       wire        [`DW-1:0]       gather_data_i_2_1,
    input       wire                        gather_valid_i_2_1,
    output      wire                        gather_ready_o_2_1,

    output      wire        [`DW-1:0]       gather_data_o_2_1,
    output      wire                        gather_valid_o_2_1,
    input       wire                        gather_ready_i_2_1,
    input       wire        [`DW-1:0]       gather_data_i_2_2,
    input       wire                        gather_valid_i_2_2,
    output      wire                        gather_ready_o_2_2,

    output      wire        [`DW-1:0]       gather_data_o_2_2,
    output      wire                        gather_valid_o_2_2,
    input       wire                        gather_ready_i_2_2,
    input       wire        [`DW-1:0]       gather_data_i_2_3,
    input       wire                        gather_valid_i_2_3,
    output      wire                        gather_ready_o_2_3,

    output      wire        [`DW-1:0]       gather_data_o_2_3,
    output      wire                        gather_valid_o_2_3,
    input       wire                        gather_ready_i_2_3,
    input       wire        [`DW-1:0]       gather_data_i_2_4,
    input       wire                        gather_valid_i_2_4,
    output      wire                        gather_ready_o_2_4,

    output      wire        [`DW-1:0]       gather_data_o_2_4,
    output      wire                        gather_valid_o_2_4,
    input       wire                        gather_ready_i_2_4,
    input       wire        [`DW-1:0]       gather_data_i_2_5,
    input       wire                        gather_valid_i_2_5,
    output      wire                        gather_ready_o_2_5,

    output      wire        [`DW-1:0]       gather_data_o_2_5,
    output      wire                        gather_valid_o_2_5,
    input       wire                        gather_ready_i_2_5,
    input       wire        [`DW-1:0]       gather_data_i_2_6,
    input       wire                        gather_valid_i_2_6,
    output      wire                        gather_ready_o_2_6,

    output      wire        [`DW-1:0]       gather_data_o_2_6,
    output      wire                        gather_valid_o_2_6,
    input       wire                        gather_ready_i_2_6,
    input       wire        [`DW-1:0]       gather_data_i_2_7,
    input       wire                        gather_valid_i_2_7,
    output      wire                        gather_ready_o_2_7,

    output      wire        [`DW-1:0]       gather_data_o_2_7,
    output      wire                        gather_valid_o_2_7,
    input       wire                        gather_ready_i_2_7,
    input       wire        [`DW-1:0]       gather_data_i_2_8,
    input       wire                        gather_valid_i_2_8,
    output      wire                        gather_ready_o_2_8,

    output      wire        [`DW-1:0]       gather_data_o_2_8,
    output      wire                        gather_valid_o_2_8,
    input       wire                        gather_ready_i_2_8,
    input       wire        [`DW-1:0]       gather_data_i_2_9,
    input       wire                        gather_valid_i_2_9,
    output      wire                        gather_ready_o_2_9,

    output      wire        [`DW-1:0]       gather_data_o_2_9,
    output      wire                        gather_valid_o_2_9,
    input       wire                        gather_ready_i_2_9,
    input       wire        [`DW-1:0]       gather_data_i_3_0,
    input       wire                        gather_valid_i_3_0,
    output      wire                        gather_ready_o_3_0,

    output      wire        [`DW-1:0]       gather_data_o_3_0,
    output      wire                        gather_valid_o_3_0,
    input       wire                        gather_ready_i_3_0,
    input       wire        [`DW-1:0]       gather_data_i_3_1,
    input       wire                        gather_valid_i_3_1,
    output      wire                        gather_ready_o_3_1,

    output      wire        [`DW-1:0]       gather_data_o_3_1,
    output      wire                        gather_valid_o_3_1,
    input       wire                        gather_ready_i_3_1,
    input       wire        [`DW-1:0]       gather_data_i_3_2,
    input       wire                        gather_valid_i_3_2,
    output      wire                        gather_ready_o_3_2,

    output      wire        [`DW-1:0]       gather_data_o_3_2,
    output      wire                        gather_valid_o_3_2,
    input       wire                        gather_ready_i_3_2,
    input       wire        [`DW-1:0]       gather_data_i_3_3,
    input       wire                        gather_valid_i_3_3,
    output      wire                        gather_ready_o_3_3,

    output      wire        [`DW-1:0]       gather_data_o_3_3,
    output      wire                        gather_valid_o_3_3,
    input       wire                        gather_ready_i_3_3,
    input       wire        [`DW-1:0]       gather_data_i_3_4,
    input       wire                        gather_valid_i_3_4,
    output      wire                        gather_ready_o_3_4,

    output      wire        [`DW-1:0]       gather_data_o_3_4,
    output      wire                        gather_valid_o_3_4,
    input       wire                        gather_ready_i_3_4,
    input       wire        [`DW-1:0]       gather_data_i_3_5,
    input       wire                        gather_valid_i_3_5,
    output      wire                        gather_ready_o_3_5,

    output      wire        [`DW-1:0]       gather_data_o_3_5,
    output      wire                        gather_valid_o_3_5,
    input       wire                        gather_ready_i_3_5,
    input       wire        [`DW-1:0]       gather_data_i_3_6,
    input       wire                        gather_valid_i_3_6,
    output      wire                        gather_ready_o_3_6,

    output      wire        [`DW-1:0]       gather_data_o_3_6,
    output      wire                        gather_valid_o_3_6,
    input       wire                        gather_ready_i_3_6,
    input       wire        [`DW-1:0]       gather_data_i_3_7,
    input       wire                        gather_valid_i_3_7,
    output      wire                        gather_ready_o_3_7,

    output      wire        [`DW-1:0]       gather_data_o_3_7,
    output      wire                        gather_valid_o_3_7,
    input       wire                        gather_ready_i_3_7,
    input       wire        [`DW-1:0]       gather_data_i_3_8,
    input       wire                        gather_valid_i_3_8,
    output      wire                        gather_ready_o_3_8,

    output      wire        [`DW-1:0]       gather_data_o_3_8,
    output      wire                        gather_valid_o_3_8,
    input       wire                        gather_ready_i_3_8,
    input       wire        [`DW-1:0]       gather_data_i_3_9,
    input       wire                        gather_valid_i_3_9,
    output      wire                        gather_ready_o_3_9,

    output      wire        [`DW-1:0]       gather_data_o_3_9,
    output      wire                        gather_valid_o_3_9,
    input       wire                        gather_ready_i_3_9,
    input       wire        [`DW-1:0]       gather_data_i_4_0,
    input       wire                        gather_valid_i_4_0,
    output      wire                        gather_ready_o_4_0,

    output      wire        [`DW-1:0]       gather_data_o_4_0,
    output      wire                        gather_valid_o_4_0,
    input       wire                        gather_ready_i_4_0,
    input       wire        [`DW-1:0]       gather_data_i_4_1,
    input       wire                        gather_valid_i_4_1,
    output      wire                        gather_ready_o_4_1,

    output      wire        [`DW-1:0]       gather_data_o_4_1,
    output      wire                        gather_valid_o_4_1,
    input       wire                        gather_ready_i_4_1,
    input       wire        [`DW-1:0]       gather_data_i_4_2,
    input       wire                        gather_valid_i_4_2,
    output      wire                        gather_ready_o_4_2,

    output      wire        [`DW-1:0]       gather_data_o_4_2,
    output      wire                        gather_valid_o_4_2,
    input       wire                        gather_ready_i_4_2,
    input       wire        [`DW-1:0]       gather_data_i_4_3,
    input       wire                        gather_valid_i_4_3,
    output      wire                        gather_ready_o_4_3,

    output      wire        [`DW-1:0]       gather_data_o_4_3,
    output      wire                        gather_valid_o_4_3,
    input       wire                        gather_ready_i_4_3,
    input       wire        [`DW-1:0]       gather_data_i_4_4,
    input       wire                        gather_valid_i_4_4,
    output      wire                        gather_ready_o_4_4,

    output      wire        [`DW-1:0]       gather_data_o_4_4,
    output      wire                        gather_valid_o_4_4,
    input       wire                        gather_ready_i_4_4,
    input       wire        [`DW-1:0]       gather_data_i_4_5,
    input       wire                        gather_valid_i_4_5,
    output      wire                        gather_ready_o_4_5,

    output      wire        [`DW-1:0]       gather_data_o_4_5,
    output      wire                        gather_valid_o_4_5,
    input       wire                        gather_ready_i_4_5,
    input       wire        [`DW-1:0]       gather_data_i_4_6,
    input       wire                        gather_valid_i_4_6,
    output      wire                        gather_ready_o_4_6,

    output      wire        [`DW-1:0]       gather_data_o_4_6,
    output      wire                        gather_valid_o_4_6,
    input       wire                        gather_ready_i_4_6,
    input       wire        [`DW-1:0]       gather_data_i_4_7,
    input       wire                        gather_valid_i_4_7,
    output      wire                        gather_ready_o_4_7,

    output      wire        [`DW-1:0]       gather_data_o_4_7,
    output      wire                        gather_valid_o_4_7,
    input       wire                        gather_ready_i_4_7,
    input       wire        [`DW-1:0]       gather_data_i_4_8,
    input       wire                        gather_valid_i_4_8,
    output      wire                        gather_ready_o_4_8,

    output      wire        [`DW-1:0]       gather_data_o_4_8,
    output      wire                        gather_valid_o_4_8,
    input       wire                        gather_ready_i_4_8,
    input       wire        [`DW-1:0]       gather_data_i_4_9,
    input       wire                        gather_valid_i_4_9,
    output      wire                        gather_ready_o_4_9,

    output      wire        [`DW-1:0]       gather_data_o_4_9,
    output      wire                        gather_valid_o_4_9,
    input       wire                        gather_ready_i_4_9
);
wire [`DW-1:0] data_stab;
wire valid_stab, ready_stab;

wire [`DW-1:0] data_flee0;
wire valid_flee0, ready_flee0;

wire [`DW-1:0] data_flee1;
wire valid_flee1, ready_flee1;

wire [`DW-1:0] data_i_cast_nw[`NOC_WIDTH][`NOC_HEIGHT], data_o_cast_nw[`NOC_WIDTH][`NOC_HEIGHT], data_i_merge_nw[`NOC_WIDTH][`NOC_HEIGHT], data_o_merge_nw[`NOC_WIDTH][`NOC_HEIGHT], data_i_gather_nw[`NOC_WIDTH][`NOC_HEIGHT], data_o_gather_nw[`NOC_WIDTH][`NOC_HEIGHT];
wire valid_i_cast_nw[`NOC_WIDTH][`NOC_HEIGHT], valid_o_cast_nw[`NOC_WIDTH][`NOC_HEIGHT], valid_i_merge_nw[`NOC_WIDTH][`NOC_HEIGHT], valid_o_merge_nw[`NOC_WIDTH][`NOC_HEIGHT], valid_i_gather_nw[`NOC_WIDTH][`NOC_HEIGHT], valid_o_gather_nw[`NOC_WIDTH][`NOC_HEIGHT];
wire ready_i_cast_nw[`NOC_WIDTH][`NOC_HEIGHT], ready_o_cast_nw[`NOC_WIDTH][`NOC_HEIGHT], ready_i_merge_nw[`NOC_WIDTH][`NOC_HEIGHT], ready_o_merge_nw[`NOC_WIDTH][`NOC_HEIGHT], ready_i_gather_nw[`NOC_WIDTH][`NOC_HEIGHT], ready_o_gather_nw[`NOC_WIDTH][`NOC_HEIGHT];

wire credit_upd[`NOC_WIDTH][`NOC_HEIGHT];

// from stab port to network
converter #(
    .out                            (1),
    .sid                            (1023)
)converter_stab(
    .clk                            (clk),
    .rstn                           (rstn),
    .valid_i_pe                     (valid_i_stab),
    .data_i_pe                      (data_i_stab),
    .ready_o_pe                     (ready_o_stab),
    .valid_o_pe                     (),
    .data_o_pe                      (),
    .ready_i_pe                     (1'b0),
    .valid_i_nw                     (1'b0),
    .data_i_nw                      ({(`DW){1'b0}}),
    .ready_o_nw                     (),
    .valid_o_nw                     (valid_stab),
    .data_o_nw                      (data_stab),
    .ready_i_nw                     (ready_stab)
);

// from flee0 port to outside
converter #(
    .out                            (0),
    .sid                            (1022)
)converter_flee0(
    .clk                            (clk),
    .rstn                           (rstn),
    .valid_i_pe                     (1'b0),
    .data_i_pe                      ({(`DW){1'b0}}),
    .ready_o_pe                     (),
    .valid_o_pe                     (valid_o_flee0),
    .data_o_pe                      (data_o_flee0),
    .ready_i_pe                     (ready_i_flee0),
    .valid_i_nw                     (valid_flee0),
    .data_i_nw                      (data_flee0),
    .ready_o_nw                     (ready_flee0),
    .valid_o_nw                     (),
    .data_o_nw                      (),
    .ready_i_nw                     (1'b0)
);

// from flee1 port to outside
converter #(
    .out                            (0),
    .sid                            (1022)
)converter_flee1(
    .clk                            (clk),
    .rstn                           (rstn),
    .valid_i_pe                     (1'b0),
    .data_i_pe                      ({(`DW){1'b0}}),
    .ready_o_pe                     (),
    .valid_o_pe                     (valid_o_flee1),
    .data_o_pe                      (data_o_flee1),
    .ready_i_pe                     (ready_i_flee1),
    .valid_i_nw                     (valid_flee1),
    .data_i_nw                      (data_flee1),
    .ready_o_nw                     (ready_flee1),
    .valid_o_nw                     (),
    .data_o_nw                      (),
    .ready_i_nw                     (1'b0)
);

cast_network cast_nw(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_cast_nw),
    .valid_i                        (valid_i_cast_nw),
    .ready_o                        (ready_o_cast_nw),
    .data_o                         (data_o_cast_nw),
    .valid_o                        (valid_o_cast_nw),
    .ready_i                        (ready_i_cast_nw),
    .data_i_stab                    (data_stab),
    .valid_i_stab                   (valid_stab),
    .ready_o_stab                   (ready_stab),
    .data_o_flee0                   (data_flee0),
    .valid_o_flee0                  (valid_flee0),
    .ready_i_flee0                  (ready_flee0),
    .data_o_flee1                   (data_flee1),
    .valid_o_flee1                  (valid_flee1),
    .ready_i_flee1                  (ready_flee1),
    .credit_upd                     (credit_upd)
);                 

merge_network merge_nw(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_merge_nw),
    .valid_i                        (valid_i_merge_nw),
    .ready_o                        (ready_o_merge_nw),
    .data_o                         (data_o_merge_nw),
    .valid_o                        (valid_o_merge_nw),
    .ready_i                        (ready_i_merge_nw)
);

gather_network gather_nw(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_gather_nw),
    .valid_i                        (valid_i_gather_nw),
    .ready_o                        (ready_o_gather_nw),
    .data_o                         (data_o_gather_nw),
    .valid_o                        (valid_o_gather_nw),
    .ready_i                        (ready_i_gather_nw)
);


network_interface #(
    .cast_out                       (cast_out_0_0),
    .gather_out                     (gather_out_0_0),
    .cast_sid                       (cast_sid_0_0),
    .gather_sid                     (gather_sid_0_0)
)ni_0_0(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[0][0]),
    .data_i_cast_nw                 (data_o_cast_nw[0][0]),
    .ready_o_cast_nw                (ready_i_cast_nw[0][0]),
    .valid_o_cast_nw                (valid_i_cast_nw[0][0]),
    .data_o_cast_nw                 (data_i_cast_nw[0][0]),
    .ready_i_cast_nw                (ready_o_cast_nw[0][0]),

    .valid_i_gather_nw              (valid_o_gather_nw[0][0]),
    .data_i_gather_nw               (data_o_gather_nw[0][0]),
    .ready_o_gather_nw              (ready_i_gather_nw[0][0]),
    .valid_o_gather_nw              (valid_i_gather_nw[0][0]),
    .data_o_gather_nw               (data_i_gather_nw[0][0]),
    .ready_i_gather_nw              (ready_o_gather_nw[0][0]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[0][0]),
    .data_i_merge_nw                (data_o_merge_nw[0][0]),
    .ready_o_merge_nw               (ready_i_merge_nw[0][0]),
    .valid_o_merge_nw               (valid_i_merge_nw[0][0]),
    .data_o_merge_nw                (data_i_merge_nw[0][0]),
    .ready_i_merge_nw               (ready_o_merge_nw[0][0]),

    .valid_i_cast_pe                (cast_valid_i_0_0),
    .data_i_cast_pe                 (cast_data_i_0_0),
    .ready_o_cast_pe                (cast_ready_o_0_0),
    .valid_o_cast_pe                (cast_valid_o_0_0),
    .data_o_cast_pe                 (cast_data_o_0_0),
    .ready_i_cast_pe                (cast_ready_i_0_0),

    .valid_i_merge_pe               (merge_valid_i_0_0),
    .data_i_merge_pe                (merge_data_i_0_0),
    .ready_o_merge_pe               (merge_ready_o_0_0),
    .valid_o_merge_pe               (merge_valid_o_0_0),
    .data_o_merge_pe                (merge_data_o_0_0),
    .ready_i_merge_pe               (merge_ready_i_0_0),

    .valid_i_gather_pe              (gather_valid_i_0_0),
    .data_i_gather_pe               (gather_data_i_0_0),
    .ready_o_gather_pe              (gather_ready_o_0_0),
    .valid_o_gather_pe              (gather_valid_o_0_0),
    .data_o_gather_pe               (gather_data_o_0_0),
    .ready_i_gather_pe              (gather_ready_i_0_0),

    .credit_upd                     (credit_upd[0][0])
);


network_interface #(
    .cast_out                       (cast_out_0_1),
    .gather_out                     (gather_out_0_1),
    .cast_sid                       (cast_sid_0_1),
    .gather_sid                     (gather_sid_0_1)
)ni_0_1(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[0][1]),
    .data_i_cast_nw                 (data_o_cast_nw[0][1]),
    .ready_o_cast_nw                (ready_i_cast_nw[0][1]),
    .valid_o_cast_nw                (valid_i_cast_nw[0][1]),
    .data_o_cast_nw                 (data_i_cast_nw[0][1]),
    .ready_i_cast_nw                (ready_o_cast_nw[0][1]),

    .valid_i_gather_nw              (valid_o_gather_nw[0][1]),
    .data_i_gather_nw               (data_o_gather_nw[0][1]),
    .ready_o_gather_nw              (ready_i_gather_nw[0][1]),
    .valid_o_gather_nw              (valid_i_gather_nw[0][1]),
    .data_o_gather_nw               (data_i_gather_nw[0][1]),
    .ready_i_gather_nw              (ready_o_gather_nw[0][1]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[0][1]),
    .data_i_merge_nw                (data_o_merge_nw[0][1]),
    .ready_o_merge_nw               (ready_i_merge_nw[0][1]),
    .valid_o_merge_nw               (valid_i_merge_nw[0][1]),
    .data_o_merge_nw                (data_i_merge_nw[0][1]),
    .ready_i_merge_nw               (ready_o_merge_nw[0][1]),

    .valid_i_cast_pe                (cast_valid_i_0_1),
    .data_i_cast_pe                 (cast_data_i_0_1),
    .ready_o_cast_pe                (cast_ready_o_0_1),
    .valid_o_cast_pe                (cast_valid_o_0_1),
    .data_o_cast_pe                 (cast_data_o_0_1),
    .ready_i_cast_pe                (cast_ready_i_0_1),

    .valid_i_merge_pe               (merge_valid_i_0_1),
    .data_i_merge_pe                (merge_data_i_0_1),
    .ready_o_merge_pe               (merge_ready_o_0_1),
    .valid_o_merge_pe               (merge_valid_o_0_1),
    .data_o_merge_pe                (merge_data_o_0_1),
    .ready_i_merge_pe               (merge_ready_i_0_1),

    .valid_i_gather_pe              (gather_valid_i_0_1),
    .data_i_gather_pe               (gather_data_i_0_1),
    .ready_o_gather_pe              (gather_ready_o_0_1),
    .valid_o_gather_pe              (gather_valid_o_0_1),
    .data_o_gather_pe               (gather_data_o_0_1),
    .ready_i_gather_pe              (gather_ready_i_0_1),

    .credit_upd                     (credit_upd[0][1])
);


network_interface #(
    .cast_out                       (cast_out_0_2),
    .gather_out                     (gather_out_0_2),
    .cast_sid                       (cast_sid_0_2),
    .gather_sid                     (gather_sid_0_2)
)ni_0_2(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[0][2]),
    .data_i_cast_nw                 (data_o_cast_nw[0][2]),
    .ready_o_cast_nw                (ready_i_cast_nw[0][2]),
    .valid_o_cast_nw                (valid_i_cast_nw[0][2]),
    .data_o_cast_nw                 (data_i_cast_nw[0][2]),
    .ready_i_cast_nw                (ready_o_cast_nw[0][2]),

    .valid_i_gather_nw              (valid_o_gather_nw[0][2]),
    .data_i_gather_nw               (data_o_gather_nw[0][2]),
    .ready_o_gather_nw              (ready_i_gather_nw[0][2]),
    .valid_o_gather_nw              (valid_i_gather_nw[0][2]),
    .data_o_gather_nw               (data_i_gather_nw[0][2]),
    .ready_i_gather_nw              (ready_o_gather_nw[0][2]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[0][2]),
    .data_i_merge_nw                (data_o_merge_nw[0][2]),
    .ready_o_merge_nw               (ready_i_merge_nw[0][2]),
    .valid_o_merge_nw               (valid_i_merge_nw[0][2]),
    .data_o_merge_nw                (data_i_merge_nw[0][2]),
    .ready_i_merge_nw               (ready_o_merge_nw[0][2]),

    .valid_i_cast_pe                (cast_valid_i_0_2),
    .data_i_cast_pe                 (cast_data_i_0_2),
    .ready_o_cast_pe                (cast_ready_o_0_2),
    .valid_o_cast_pe                (cast_valid_o_0_2),
    .data_o_cast_pe                 (cast_data_o_0_2),
    .ready_i_cast_pe                (cast_ready_i_0_2),

    .valid_i_merge_pe               (merge_valid_i_0_2),
    .data_i_merge_pe                (merge_data_i_0_2),
    .ready_o_merge_pe               (merge_ready_o_0_2),
    .valid_o_merge_pe               (merge_valid_o_0_2),
    .data_o_merge_pe                (merge_data_o_0_2),
    .ready_i_merge_pe               (merge_ready_i_0_2),

    .valid_i_gather_pe              (gather_valid_i_0_2),
    .data_i_gather_pe               (gather_data_i_0_2),
    .ready_o_gather_pe              (gather_ready_o_0_2),
    .valid_o_gather_pe              (gather_valid_o_0_2),
    .data_o_gather_pe               (gather_data_o_0_2),
    .ready_i_gather_pe              (gather_ready_i_0_2),

    .credit_upd                     (credit_upd[0][2])
);


network_interface #(
    .cast_out                       (cast_out_0_3),
    .gather_out                     (gather_out_0_3),
    .cast_sid                       (cast_sid_0_3),
    .gather_sid                     (gather_sid_0_3)
)ni_0_3(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[0][3]),
    .data_i_cast_nw                 (data_o_cast_nw[0][3]),
    .ready_o_cast_nw                (ready_i_cast_nw[0][3]),
    .valid_o_cast_nw                (valid_i_cast_nw[0][3]),
    .data_o_cast_nw                 (data_i_cast_nw[0][3]),
    .ready_i_cast_nw                (ready_o_cast_nw[0][3]),

    .valid_i_gather_nw              (valid_o_gather_nw[0][3]),
    .data_i_gather_nw               (data_o_gather_nw[0][3]),
    .ready_o_gather_nw              (ready_i_gather_nw[0][3]),
    .valid_o_gather_nw              (valid_i_gather_nw[0][3]),
    .data_o_gather_nw               (data_i_gather_nw[0][3]),
    .ready_i_gather_nw              (ready_o_gather_nw[0][3]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[0][3]),
    .data_i_merge_nw                (data_o_merge_nw[0][3]),
    .ready_o_merge_nw               (ready_i_merge_nw[0][3]),
    .valid_o_merge_nw               (valid_i_merge_nw[0][3]),
    .data_o_merge_nw                (data_i_merge_nw[0][3]),
    .ready_i_merge_nw               (ready_o_merge_nw[0][3]),

    .valid_i_cast_pe                (cast_valid_i_0_3),
    .data_i_cast_pe                 (cast_data_i_0_3),
    .ready_o_cast_pe                (cast_ready_o_0_3),
    .valid_o_cast_pe                (cast_valid_o_0_3),
    .data_o_cast_pe                 (cast_data_o_0_3),
    .ready_i_cast_pe                (cast_ready_i_0_3),

    .valid_i_merge_pe               (merge_valid_i_0_3),
    .data_i_merge_pe                (merge_data_i_0_3),
    .ready_o_merge_pe               (merge_ready_o_0_3),
    .valid_o_merge_pe               (merge_valid_o_0_3),
    .data_o_merge_pe                (merge_data_o_0_3),
    .ready_i_merge_pe               (merge_ready_i_0_3),

    .valid_i_gather_pe              (gather_valid_i_0_3),
    .data_i_gather_pe               (gather_data_i_0_3),
    .ready_o_gather_pe              (gather_ready_o_0_3),
    .valid_o_gather_pe              (gather_valid_o_0_3),
    .data_o_gather_pe               (gather_data_o_0_3),
    .ready_i_gather_pe              (gather_ready_i_0_3),

    .credit_upd                     (credit_upd[0][3])
);


network_interface #(
    .cast_out                       (cast_out_0_4),
    .gather_out                     (gather_out_0_4),
    .cast_sid                       (cast_sid_0_4),
    .gather_sid                     (gather_sid_0_4)
)ni_0_4(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[0][4]),
    .data_i_cast_nw                 (data_o_cast_nw[0][4]),
    .ready_o_cast_nw                (ready_i_cast_nw[0][4]),
    .valid_o_cast_nw                (valid_i_cast_nw[0][4]),
    .data_o_cast_nw                 (data_i_cast_nw[0][4]),
    .ready_i_cast_nw                (ready_o_cast_nw[0][4]),

    .valid_i_gather_nw              (valid_o_gather_nw[0][4]),
    .data_i_gather_nw               (data_o_gather_nw[0][4]),
    .ready_o_gather_nw              (ready_i_gather_nw[0][4]),
    .valid_o_gather_nw              (valid_i_gather_nw[0][4]),
    .data_o_gather_nw               (data_i_gather_nw[0][4]),
    .ready_i_gather_nw              (ready_o_gather_nw[0][4]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[0][4]),
    .data_i_merge_nw                (data_o_merge_nw[0][4]),
    .ready_o_merge_nw               (ready_i_merge_nw[0][4]),
    .valid_o_merge_nw               (valid_i_merge_nw[0][4]),
    .data_o_merge_nw                (data_i_merge_nw[0][4]),
    .ready_i_merge_nw               (ready_o_merge_nw[0][4]),

    .valid_i_cast_pe                (cast_valid_i_0_4),
    .data_i_cast_pe                 (cast_data_i_0_4),
    .ready_o_cast_pe                (cast_ready_o_0_4),
    .valid_o_cast_pe                (cast_valid_o_0_4),
    .data_o_cast_pe                 (cast_data_o_0_4),
    .ready_i_cast_pe                (cast_ready_i_0_4),

    .valid_i_merge_pe               (merge_valid_i_0_4),
    .data_i_merge_pe                (merge_data_i_0_4),
    .ready_o_merge_pe               (merge_ready_o_0_4),
    .valid_o_merge_pe               (merge_valid_o_0_4),
    .data_o_merge_pe                (merge_data_o_0_4),
    .ready_i_merge_pe               (merge_ready_i_0_4),

    .valid_i_gather_pe              (gather_valid_i_0_4),
    .data_i_gather_pe               (gather_data_i_0_4),
    .ready_o_gather_pe              (gather_ready_o_0_4),
    .valid_o_gather_pe              (gather_valid_o_0_4),
    .data_o_gather_pe               (gather_data_o_0_4),
    .ready_i_gather_pe              (gather_ready_i_0_4),

    .credit_upd                     (credit_upd[0][4])
);


network_interface #(
    .cast_out                       (cast_out_0_5),
    .gather_out                     (gather_out_0_5),
    .cast_sid                       (cast_sid_0_5),
    .gather_sid                     (gather_sid_0_5)
)ni_0_5(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[0][5]),
    .data_i_cast_nw                 (data_o_cast_nw[0][5]),
    .ready_o_cast_nw                (ready_i_cast_nw[0][5]),
    .valid_o_cast_nw                (valid_i_cast_nw[0][5]),
    .data_o_cast_nw                 (data_i_cast_nw[0][5]),
    .ready_i_cast_nw                (ready_o_cast_nw[0][5]),

    .valid_i_gather_nw              (valid_o_gather_nw[0][5]),
    .data_i_gather_nw               (data_o_gather_nw[0][5]),
    .ready_o_gather_nw              (ready_i_gather_nw[0][5]),
    .valid_o_gather_nw              (valid_i_gather_nw[0][5]),
    .data_o_gather_nw               (data_i_gather_nw[0][5]),
    .ready_i_gather_nw              (ready_o_gather_nw[0][5]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[0][5]),
    .data_i_merge_nw                (data_o_merge_nw[0][5]),
    .ready_o_merge_nw               (ready_i_merge_nw[0][5]),
    .valid_o_merge_nw               (valid_i_merge_nw[0][5]),
    .data_o_merge_nw                (data_i_merge_nw[0][5]),
    .ready_i_merge_nw               (ready_o_merge_nw[0][5]),

    .valid_i_cast_pe                (cast_valid_i_0_5),
    .data_i_cast_pe                 (cast_data_i_0_5),
    .ready_o_cast_pe                (cast_ready_o_0_5),
    .valid_o_cast_pe                (cast_valid_o_0_5),
    .data_o_cast_pe                 (cast_data_o_0_5),
    .ready_i_cast_pe                (cast_ready_i_0_5),

    .valid_i_merge_pe               (merge_valid_i_0_5),
    .data_i_merge_pe                (merge_data_i_0_5),
    .ready_o_merge_pe               (merge_ready_o_0_5),
    .valid_o_merge_pe               (merge_valid_o_0_5),
    .data_o_merge_pe                (merge_data_o_0_5),
    .ready_i_merge_pe               (merge_ready_i_0_5),

    .valid_i_gather_pe              (gather_valid_i_0_5),
    .data_i_gather_pe               (gather_data_i_0_5),
    .ready_o_gather_pe              (gather_ready_o_0_5),
    .valid_o_gather_pe              (gather_valid_o_0_5),
    .data_o_gather_pe               (gather_data_o_0_5),
    .ready_i_gather_pe              (gather_ready_i_0_5),

    .credit_upd                     (credit_upd[0][5])
);


network_interface #(
    .cast_out                       (cast_out_0_6),
    .gather_out                     (gather_out_0_6),
    .cast_sid                       (cast_sid_0_6),
    .gather_sid                     (gather_sid_0_6)
)ni_0_6(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[0][6]),
    .data_i_cast_nw                 (data_o_cast_nw[0][6]),
    .ready_o_cast_nw                (ready_i_cast_nw[0][6]),
    .valid_o_cast_nw                (valid_i_cast_nw[0][6]),
    .data_o_cast_nw                 (data_i_cast_nw[0][6]),
    .ready_i_cast_nw                (ready_o_cast_nw[0][6]),

    .valid_i_gather_nw              (valid_o_gather_nw[0][6]),
    .data_i_gather_nw               (data_o_gather_nw[0][6]),
    .ready_o_gather_nw              (ready_i_gather_nw[0][6]),
    .valid_o_gather_nw              (valid_i_gather_nw[0][6]),
    .data_o_gather_nw               (data_i_gather_nw[0][6]),
    .ready_i_gather_nw              (ready_o_gather_nw[0][6]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[0][6]),
    .data_i_merge_nw                (data_o_merge_nw[0][6]),
    .ready_o_merge_nw               (ready_i_merge_nw[0][6]),
    .valid_o_merge_nw               (valid_i_merge_nw[0][6]),
    .data_o_merge_nw                (data_i_merge_nw[0][6]),
    .ready_i_merge_nw               (ready_o_merge_nw[0][6]),

    .valid_i_cast_pe                (cast_valid_i_0_6),
    .data_i_cast_pe                 (cast_data_i_0_6),
    .ready_o_cast_pe                (cast_ready_o_0_6),
    .valid_o_cast_pe                (cast_valid_o_0_6),
    .data_o_cast_pe                 (cast_data_o_0_6),
    .ready_i_cast_pe                (cast_ready_i_0_6),

    .valid_i_merge_pe               (merge_valid_i_0_6),
    .data_i_merge_pe                (merge_data_i_0_6),
    .ready_o_merge_pe               (merge_ready_o_0_6),
    .valid_o_merge_pe               (merge_valid_o_0_6),
    .data_o_merge_pe                (merge_data_o_0_6),
    .ready_i_merge_pe               (merge_ready_i_0_6),

    .valid_i_gather_pe              (gather_valid_i_0_6),
    .data_i_gather_pe               (gather_data_i_0_6),
    .ready_o_gather_pe              (gather_ready_o_0_6),
    .valid_o_gather_pe              (gather_valid_o_0_6),
    .data_o_gather_pe               (gather_data_o_0_6),
    .ready_i_gather_pe              (gather_ready_i_0_6),

    .credit_upd                     (credit_upd[0][6])
);


network_interface #(
    .cast_out                       (cast_out_0_7),
    .gather_out                     (gather_out_0_7),
    .cast_sid                       (cast_sid_0_7),
    .gather_sid                     (gather_sid_0_7)
)ni_0_7(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[0][7]),
    .data_i_cast_nw                 (data_o_cast_nw[0][7]),
    .ready_o_cast_nw                (ready_i_cast_nw[0][7]),
    .valid_o_cast_nw                (valid_i_cast_nw[0][7]),
    .data_o_cast_nw                 (data_i_cast_nw[0][7]),
    .ready_i_cast_nw                (ready_o_cast_nw[0][7]),

    .valid_i_gather_nw              (valid_o_gather_nw[0][7]),
    .data_i_gather_nw               (data_o_gather_nw[0][7]),
    .ready_o_gather_nw              (ready_i_gather_nw[0][7]),
    .valid_o_gather_nw              (valid_i_gather_nw[0][7]),
    .data_o_gather_nw               (data_i_gather_nw[0][7]),
    .ready_i_gather_nw              (ready_o_gather_nw[0][7]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[0][7]),
    .data_i_merge_nw                (data_o_merge_nw[0][7]),
    .ready_o_merge_nw               (ready_i_merge_nw[0][7]),
    .valid_o_merge_nw               (valid_i_merge_nw[0][7]),
    .data_o_merge_nw                (data_i_merge_nw[0][7]),
    .ready_i_merge_nw               (ready_o_merge_nw[0][7]),

    .valid_i_cast_pe                (cast_valid_i_0_7),
    .data_i_cast_pe                 (cast_data_i_0_7),
    .ready_o_cast_pe                (cast_ready_o_0_7),
    .valid_o_cast_pe                (cast_valid_o_0_7),
    .data_o_cast_pe                 (cast_data_o_0_7),
    .ready_i_cast_pe                (cast_ready_i_0_7),

    .valid_i_merge_pe               (merge_valid_i_0_7),
    .data_i_merge_pe                (merge_data_i_0_7),
    .ready_o_merge_pe               (merge_ready_o_0_7),
    .valid_o_merge_pe               (merge_valid_o_0_7),
    .data_o_merge_pe                (merge_data_o_0_7),
    .ready_i_merge_pe               (merge_ready_i_0_7),

    .valid_i_gather_pe              (gather_valid_i_0_7),
    .data_i_gather_pe               (gather_data_i_0_7),
    .ready_o_gather_pe              (gather_ready_o_0_7),
    .valid_o_gather_pe              (gather_valid_o_0_7),
    .data_o_gather_pe               (gather_data_o_0_7),
    .ready_i_gather_pe              (gather_ready_i_0_7),

    .credit_upd                     (credit_upd[0][7])
);


network_interface #(
    .cast_out                       (cast_out_0_8),
    .gather_out                     (gather_out_0_8),
    .cast_sid                       (cast_sid_0_8),
    .gather_sid                     (gather_sid_0_8)
)ni_0_8(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[0][8]),
    .data_i_cast_nw                 (data_o_cast_nw[0][8]),
    .ready_o_cast_nw                (ready_i_cast_nw[0][8]),
    .valid_o_cast_nw                (valid_i_cast_nw[0][8]),
    .data_o_cast_nw                 (data_i_cast_nw[0][8]),
    .ready_i_cast_nw                (ready_o_cast_nw[0][8]),

    .valid_i_gather_nw              (valid_o_gather_nw[0][8]),
    .data_i_gather_nw               (data_o_gather_nw[0][8]),
    .ready_o_gather_nw              (ready_i_gather_nw[0][8]),
    .valid_o_gather_nw              (valid_i_gather_nw[0][8]),
    .data_o_gather_nw               (data_i_gather_nw[0][8]),
    .ready_i_gather_nw              (ready_o_gather_nw[0][8]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[0][8]),
    .data_i_merge_nw                (data_o_merge_nw[0][8]),
    .ready_o_merge_nw               (ready_i_merge_nw[0][8]),
    .valid_o_merge_nw               (valid_i_merge_nw[0][8]),
    .data_o_merge_nw                (data_i_merge_nw[0][8]),
    .ready_i_merge_nw               (ready_o_merge_nw[0][8]),

    .valid_i_cast_pe                (cast_valid_i_0_8),
    .data_i_cast_pe                 (cast_data_i_0_8),
    .ready_o_cast_pe                (cast_ready_o_0_8),
    .valid_o_cast_pe                (cast_valid_o_0_8),
    .data_o_cast_pe                 (cast_data_o_0_8),
    .ready_i_cast_pe                (cast_ready_i_0_8),

    .valid_i_merge_pe               (merge_valid_i_0_8),
    .data_i_merge_pe                (merge_data_i_0_8),
    .ready_o_merge_pe               (merge_ready_o_0_8),
    .valid_o_merge_pe               (merge_valid_o_0_8),
    .data_o_merge_pe                (merge_data_o_0_8),
    .ready_i_merge_pe               (merge_ready_i_0_8),

    .valid_i_gather_pe              (gather_valid_i_0_8),
    .data_i_gather_pe               (gather_data_i_0_8),
    .ready_o_gather_pe              (gather_ready_o_0_8),
    .valid_o_gather_pe              (gather_valid_o_0_8),
    .data_o_gather_pe               (gather_data_o_0_8),
    .ready_i_gather_pe              (gather_ready_i_0_8),

    .credit_upd                     (credit_upd[0][8])
);


network_interface #(
    .cast_out                       (cast_out_0_9),
    .gather_out                     (gather_out_0_9),
    .cast_sid                       (cast_sid_0_9),
    .gather_sid                     (gather_sid_0_9)
)ni_0_9(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[0][9]),
    .data_i_cast_nw                 (data_o_cast_nw[0][9]),
    .ready_o_cast_nw                (ready_i_cast_nw[0][9]),
    .valid_o_cast_nw                (valid_i_cast_nw[0][9]),
    .data_o_cast_nw                 (data_i_cast_nw[0][9]),
    .ready_i_cast_nw                (ready_o_cast_nw[0][9]),

    .valid_i_gather_nw              (valid_o_gather_nw[0][9]),
    .data_i_gather_nw               (data_o_gather_nw[0][9]),
    .ready_o_gather_nw              (ready_i_gather_nw[0][9]),
    .valid_o_gather_nw              (valid_i_gather_nw[0][9]),
    .data_o_gather_nw               (data_i_gather_nw[0][9]),
    .ready_i_gather_nw              (ready_o_gather_nw[0][9]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[0][9]),
    .data_i_merge_nw                (data_o_merge_nw[0][9]),
    .ready_o_merge_nw               (ready_i_merge_nw[0][9]),
    .valid_o_merge_nw               (valid_i_merge_nw[0][9]),
    .data_o_merge_nw                (data_i_merge_nw[0][9]),
    .ready_i_merge_nw               (ready_o_merge_nw[0][9]),

    .valid_i_cast_pe                (cast_valid_i_0_9),
    .data_i_cast_pe                 (cast_data_i_0_9),
    .ready_o_cast_pe                (cast_ready_o_0_9),
    .valid_o_cast_pe                (cast_valid_o_0_9),
    .data_o_cast_pe                 (cast_data_o_0_9),
    .ready_i_cast_pe                (cast_ready_i_0_9),

    .valid_i_merge_pe               (merge_valid_i_0_9),
    .data_i_merge_pe                (merge_data_i_0_9),
    .ready_o_merge_pe               (merge_ready_o_0_9),
    .valid_o_merge_pe               (merge_valid_o_0_9),
    .data_o_merge_pe                (merge_data_o_0_9),
    .ready_i_merge_pe               (merge_ready_i_0_9),

    .valid_i_gather_pe              (gather_valid_i_0_9),
    .data_i_gather_pe               (gather_data_i_0_9),
    .ready_o_gather_pe              (gather_ready_o_0_9),
    .valid_o_gather_pe              (gather_valid_o_0_9),
    .data_o_gather_pe               (gather_data_o_0_9),
    .ready_i_gather_pe              (gather_ready_i_0_9),

    .credit_upd                     (credit_upd[0][9])
);


network_interface #(
    .cast_out                       (cast_out_1_0),
    .gather_out                     (gather_out_1_0),
    .cast_sid                       (cast_sid_1_0),
    .gather_sid                     (gather_sid_1_0)
)ni_1_0(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[1][0]),
    .data_i_cast_nw                 (data_o_cast_nw[1][0]),
    .ready_o_cast_nw                (ready_i_cast_nw[1][0]),
    .valid_o_cast_nw                (valid_i_cast_nw[1][0]),
    .data_o_cast_nw                 (data_i_cast_nw[1][0]),
    .ready_i_cast_nw                (ready_o_cast_nw[1][0]),

    .valid_i_gather_nw              (valid_o_gather_nw[1][0]),
    .data_i_gather_nw               (data_o_gather_nw[1][0]),
    .ready_o_gather_nw              (ready_i_gather_nw[1][0]),
    .valid_o_gather_nw              (valid_i_gather_nw[1][0]),
    .data_o_gather_nw               (data_i_gather_nw[1][0]),
    .ready_i_gather_nw              (ready_o_gather_nw[1][0]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[1][0]),
    .data_i_merge_nw                (data_o_merge_nw[1][0]),
    .ready_o_merge_nw               (ready_i_merge_nw[1][0]),
    .valid_o_merge_nw               (valid_i_merge_nw[1][0]),
    .data_o_merge_nw                (data_i_merge_nw[1][0]),
    .ready_i_merge_nw               (ready_o_merge_nw[1][0]),

    .valid_i_cast_pe                (cast_valid_i_1_0),
    .data_i_cast_pe                 (cast_data_i_1_0),
    .ready_o_cast_pe                (cast_ready_o_1_0),
    .valid_o_cast_pe                (cast_valid_o_1_0),
    .data_o_cast_pe                 (cast_data_o_1_0),
    .ready_i_cast_pe                (cast_ready_i_1_0),

    .valid_i_merge_pe               (merge_valid_i_1_0),
    .data_i_merge_pe                (merge_data_i_1_0),
    .ready_o_merge_pe               (merge_ready_o_1_0),
    .valid_o_merge_pe               (merge_valid_o_1_0),
    .data_o_merge_pe                (merge_data_o_1_0),
    .ready_i_merge_pe               (merge_ready_i_1_0),

    .valid_i_gather_pe              (gather_valid_i_1_0),
    .data_i_gather_pe               (gather_data_i_1_0),
    .ready_o_gather_pe              (gather_ready_o_1_0),
    .valid_o_gather_pe              (gather_valid_o_1_0),
    .data_o_gather_pe               (gather_data_o_1_0),
    .ready_i_gather_pe              (gather_ready_i_1_0),

    .credit_upd                     (credit_upd[1][0])
);


network_interface #(
    .cast_out                       (cast_out_1_1),
    .gather_out                     (gather_out_1_1),
    .cast_sid                       (cast_sid_1_1),
    .gather_sid                     (gather_sid_1_1)
)ni_1_1(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[1][1]),
    .data_i_cast_nw                 (data_o_cast_nw[1][1]),
    .ready_o_cast_nw                (ready_i_cast_nw[1][1]),
    .valid_o_cast_nw                (valid_i_cast_nw[1][1]),
    .data_o_cast_nw                 (data_i_cast_nw[1][1]),
    .ready_i_cast_nw                (ready_o_cast_nw[1][1]),

    .valid_i_gather_nw              (valid_o_gather_nw[1][1]),
    .data_i_gather_nw               (data_o_gather_nw[1][1]),
    .ready_o_gather_nw              (ready_i_gather_nw[1][1]),
    .valid_o_gather_nw              (valid_i_gather_nw[1][1]),
    .data_o_gather_nw               (data_i_gather_nw[1][1]),
    .ready_i_gather_nw              (ready_o_gather_nw[1][1]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[1][1]),
    .data_i_merge_nw                (data_o_merge_nw[1][1]),
    .ready_o_merge_nw               (ready_i_merge_nw[1][1]),
    .valid_o_merge_nw               (valid_i_merge_nw[1][1]),
    .data_o_merge_nw                (data_i_merge_nw[1][1]),
    .ready_i_merge_nw               (ready_o_merge_nw[1][1]),

    .valid_i_cast_pe                (cast_valid_i_1_1),
    .data_i_cast_pe                 (cast_data_i_1_1),
    .ready_o_cast_pe                (cast_ready_o_1_1),
    .valid_o_cast_pe                (cast_valid_o_1_1),
    .data_o_cast_pe                 (cast_data_o_1_1),
    .ready_i_cast_pe                (cast_ready_i_1_1),

    .valid_i_merge_pe               (merge_valid_i_1_1),
    .data_i_merge_pe                (merge_data_i_1_1),
    .ready_o_merge_pe               (merge_ready_o_1_1),
    .valid_o_merge_pe               (merge_valid_o_1_1),
    .data_o_merge_pe                (merge_data_o_1_1),
    .ready_i_merge_pe               (merge_ready_i_1_1),

    .valid_i_gather_pe              (gather_valid_i_1_1),
    .data_i_gather_pe               (gather_data_i_1_1),
    .ready_o_gather_pe              (gather_ready_o_1_1),
    .valid_o_gather_pe              (gather_valid_o_1_1),
    .data_o_gather_pe               (gather_data_o_1_1),
    .ready_i_gather_pe              (gather_ready_i_1_1),

    .credit_upd                     (credit_upd[1][1])
);


network_interface #(
    .cast_out                       (cast_out_1_2),
    .gather_out                     (gather_out_1_2),
    .cast_sid                       (cast_sid_1_2),
    .gather_sid                     (gather_sid_1_2)
)ni_1_2(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[1][2]),
    .data_i_cast_nw                 (data_o_cast_nw[1][2]),
    .ready_o_cast_nw                (ready_i_cast_nw[1][2]),
    .valid_o_cast_nw                (valid_i_cast_nw[1][2]),
    .data_o_cast_nw                 (data_i_cast_nw[1][2]),
    .ready_i_cast_nw                (ready_o_cast_nw[1][2]),

    .valid_i_gather_nw              (valid_o_gather_nw[1][2]),
    .data_i_gather_nw               (data_o_gather_nw[1][2]),
    .ready_o_gather_nw              (ready_i_gather_nw[1][2]),
    .valid_o_gather_nw              (valid_i_gather_nw[1][2]),
    .data_o_gather_nw               (data_i_gather_nw[1][2]),
    .ready_i_gather_nw              (ready_o_gather_nw[1][2]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[1][2]),
    .data_i_merge_nw                (data_o_merge_nw[1][2]),
    .ready_o_merge_nw               (ready_i_merge_nw[1][2]),
    .valid_o_merge_nw               (valid_i_merge_nw[1][2]),
    .data_o_merge_nw                (data_i_merge_nw[1][2]),
    .ready_i_merge_nw               (ready_o_merge_nw[1][2]),

    .valid_i_cast_pe                (cast_valid_i_1_2),
    .data_i_cast_pe                 (cast_data_i_1_2),
    .ready_o_cast_pe                (cast_ready_o_1_2),
    .valid_o_cast_pe                (cast_valid_o_1_2),
    .data_o_cast_pe                 (cast_data_o_1_2),
    .ready_i_cast_pe                (cast_ready_i_1_2),

    .valid_i_merge_pe               (merge_valid_i_1_2),
    .data_i_merge_pe                (merge_data_i_1_2),
    .ready_o_merge_pe               (merge_ready_o_1_2),
    .valid_o_merge_pe               (merge_valid_o_1_2),
    .data_o_merge_pe                (merge_data_o_1_2),
    .ready_i_merge_pe               (merge_ready_i_1_2),

    .valid_i_gather_pe              (gather_valid_i_1_2),
    .data_i_gather_pe               (gather_data_i_1_2),
    .ready_o_gather_pe              (gather_ready_o_1_2),
    .valid_o_gather_pe              (gather_valid_o_1_2),
    .data_o_gather_pe               (gather_data_o_1_2),
    .ready_i_gather_pe              (gather_ready_i_1_2),

    .credit_upd                     (credit_upd[1][2])
);


network_interface #(
    .cast_out                       (cast_out_1_3),
    .gather_out                     (gather_out_1_3),
    .cast_sid                       (cast_sid_1_3),
    .gather_sid                     (gather_sid_1_3)
)ni_1_3(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[1][3]),
    .data_i_cast_nw                 (data_o_cast_nw[1][3]),
    .ready_o_cast_nw                (ready_i_cast_nw[1][3]),
    .valid_o_cast_nw                (valid_i_cast_nw[1][3]),
    .data_o_cast_nw                 (data_i_cast_nw[1][3]),
    .ready_i_cast_nw                (ready_o_cast_nw[1][3]),

    .valid_i_gather_nw              (valid_o_gather_nw[1][3]),
    .data_i_gather_nw               (data_o_gather_nw[1][3]),
    .ready_o_gather_nw              (ready_i_gather_nw[1][3]),
    .valid_o_gather_nw              (valid_i_gather_nw[1][3]),
    .data_o_gather_nw               (data_i_gather_nw[1][3]),
    .ready_i_gather_nw              (ready_o_gather_nw[1][3]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[1][3]),
    .data_i_merge_nw                (data_o_merge_nw[1][3]),
    .ready_o_merge_nw               (ready_i_merge_nw[1][3]),
    .valid_o_merge_nw               (valid_i_merge_nw[1][3]),
    .data_o_merge_nw                (data_i_merge_nw[1][3]),
    .ready_i_merge_nw               (ready_o_merge_nw[1][3]),

    .valid_i_cast_pe                (cast_valid_i_1_3),
    .data_i_cast_pe                 (cast_data_i_1_3),
    .ready_o_cast_pe                (cast_ready_o_1_3),
    .valid_o_cast_pe                (cast_valid_o_1_3),
    .data_o_cast_pe                 (cast_data_o_1_3),
    .ready_i_cast_pe                (cast_ready_i_1_3),

    .valid_i_merge_pe               (merge_valid_i_1_3),
    .data_i_merge_pe                (merge_data_i_1_3),
    .ready_o_merge_pe               (merge_ready_o_1_3),
    .valid_o_merge_pe               (merge_valid_o_1_3),
    .data_o_merge_pe                (merge_data_o_1_3),
    .ready_i_merge_pe               (merge_ready_i_1_3),

    .valid_i_gather_pe              (gather_valid_i_1_3),
    .data_i_gather_pe               (gather_data_i_1_3),
    .ready_o_gather_pe              (gather_ready_o_1_3),
    .valid_o_gather_pe              (gather_valid_o_1_3),
    .data_o_gather_pe               (gather_data_o_1_3),
    .ready_i_gather_pe              (gather_ready_i_1_3),

    .credit_upd                     (credit_upd[1][3])
);


network_interface #(
    .cast_out                       (cast_out_1_4),
    .gather_out                     (gather_out_1_4),
    .cast_sid                       (cast_sid_1_4),
    .gather_sid                     (gather_sid_1_4)
)ni_1_4(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[1][4]),
    .data_i_cast_nw                 (data_o_cast_nw[1][4]),
    .ready_o_cast_nw                (ready_i_cast_nw[1][4]),
    .valid_o_cast_nw                (valid_i_cast_nw[1][4]),
    .data_o_cast_nw                 (data_i_cast_nw[1][4]),
    .ready_i_cast_nw                (ready_o_cast_nw[1][4]),

    .valid_i_gather_nw              (valid_o_gather_nw[1][4]),
    .data_i_gather_nw               (data_o_gather_nw[1][4]),
    .ready_o_gather_nw              (ready_i_gather_nw[1][4]),
    .valid_o_gather_nw              (valid_i_gather_nw[1][4]),
    .data_o_gather_nw               (data_i_gather_nw[1][4]),
    .ready_i_gather_nw              (ready_o_gather_nw[1][4]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[1][4]),
    .data_i_merge_nw                (data_o_merge_nw[1][4]),
    .ready_o_merge_nw               (ready_i_merge_nw[1][4]),
    .valid_o_merge_nw               (valid_i_merge_nw[1][4]),
    .data_o_merge_nw                (data_i_merge_nw[1][4]),
    .ready_i_merge_nw               (ready_o_merge_nw[1][4]),

    .valid_i_cast_pe                (cast_valid_i_1_4),
    .data_i_cast_pe                 (cast_data_i_1_4),
    .ready_o_cast_pe                (cast_ready_o_1_4),
    .valid_o_cast_pe                (cast_valid_o_1_4),
    .data_o_cast_pe                 (cast_data_o_1_4),
    .ready_i_cast_pe                (cast_ready_i_1_4),

    .valid_i_merge_pe               (merge_valid_i_1_4),
    .data_i_merge_pe                (merge_data_i_1_4),
    .ready_o_merge_pe               (merge_ready_o_1_4),
    .valid_o_merge_pe               (merge_valid_o_1_4),
    .data_o_merge_pe                (merge_data_o_1_4),
    .ready_i_merge_pe               (merge_ready_i_1_4),

    .valid_i_gather_pe              (gather_valid_i_1_4),
    .data_i_gather_pe               (gather_data_i_1_4),
    .ready_o_gather_pe              (gather_ready_o_1_4),
    .valid_o_gather_pe              (gather_valid_o_1_4),
    .data_o_gather_pe               (gather_data_o_1_4),
    .ready_i_gather_pe              (gather_ready_i_1_4),

    .credit_upd                     (credit_upd[1][4])
);


network_interface #(
    .cast_out                       (cast_out_1_5),
    .gather_out                     (gather_out_1_5),
    .cast_sid                       (cast_sid_1_5),
    .gather_sid                     (gather_sid_1_5)
)ni_1_5(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[1][5]),
    .data_i_cast_nw                 (data_o_cast_nw[1][5]),
    .ready_o_cast_nw                (ready_i_cast_nw[1][5]),
    .valid_o_cast_nw                (valid_i_cast_nw[1][5]),
    .data_o_cast_nw                 (data_i_cast_nw[1][5]),
    .ready_i_cast_nw                (ready_o_cast_nw[1][5]),

    .valid_i_gather_nw              (valid_o_gather_nw[1][5]),
    .data_i_gather_nw               (data_o_gather_nw[1][5]),
    .ready_o_gather_nw              (ready_i_gather_nw[1][5]),
    .valid_o_gather_nw              (valid_i_gather_nw[1][5]),
    .data_o_gather_nw               (data_i_gather_nw[1][5]),
    .ready_i_gather_nw              (ready_o_gather_nw[1][5]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[1][5]),
    .data_i_merge_nw                (data_o_merge_nw[1][5]),
    .ready_o_merge_nw               (ready_i_merge_nw[1][5]),
    .valid_o_merge_nw               (valid_i_merge_nw[1][5]),
    .data_o_merge_nw                (data_i_merge_nw[1][5]),
    .ready_i_merge_nw               (ready_o_merge_nw[1][5]),

    .valid_i_cast_pe                (cast_valid_i_1_5),
    .data_i_cast_pe                 (cast_data_i_1_5),
    .ready_o_cast_pe                (cast_ready_o_1_5),
    .valid_o_cast_pe                (cast_valid_o_1_5),
    .data_o_cast_pe                 (cast_data_o_1_5),
    .ready_i_cast_pe                (cast_ready_i_1_5),

    .valid_i_merge_pe               (merge_valid_i_1_5),
    .data_i_merge_pe                (merge_data_i_1_5),
    .ready_o_merge_pe               (merge_ready_o_1_5),
    .valid_o_merge_pe               (merge_valid_o_1_5),
    .data_o_merge_pe                (merge_data_o_1_5),
    .ready_i_merge_pe               (merge_ready_i_1_5),

    .valid_i_gather_pe              (gather_valid_i_1_5),
    .data_i_gather_pe               (gather_data_i_1_5),
    .ready_o_gather_pe              (gather_ready_o_1_5),
    .valid_o_gather_pe              (gather_valid_o_1_5),
    .data_o_gather_pe               (gather_data_o_1_5),
    .ready_i_gather_pe              (gather_ready_i_1_5),

    .credit_upd                     (credit_upd[1][5])
);


network_interface #(
    .cast_out                       (cast_out_1_6),
    .gather_out                     (gather_out_1_6),
    .cast_sid                       (cast_sid_1_6),
    .gather_sid                     (gather_sid_1_6)
)ni_1_6(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[1][6]),
    .data_i_cast_nw                 (data_o_cast_nw[1][6]),
    .ready_o_cast_nw                (ready_i_cast_nw[1][6]),
    .valid_o_cast_nw                (valid_i_cast_nw[1][6]),
    .data_o_cast_nw                 (data_i_cast_nw[1][6]),
    .ready_i_cast_nw                (ready_o_cast_nw[1][6]),

    .valid_i_gather_nw              (valid_o_gather_nw[1][6]),
    .data_i_gather_nw               (data_o_gather_nw[1][6]),
    .ready_o_gather_nw              (ready_i_gather_nw[1][6]),
    .valid_o_gather_nw              (valid_i_gather_nw[1][6]),
    .data_o_gather_nw               (data_i_gather_nw[1][6]),
    .ready_i_gather_nw              (ready_o_gather_nw[1][6]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[1][6]),
    .data_i_merge_nw                (data_o_merge_nw[1][6]),
    .ready_o_merge_nw               (ready_i_merge_nw[1][6]),
    .valid_o_merge_nw               (valid_i_merge_nw[1][6]),
    .data_o_merge_nw                (data_i_merge_nw[1][6]),
    .ready_i_merge_nw               (ready_o_merge_nw[1][6]),

    .valid_i_cast_pe                (cast_valid_i_1_6),
    .data_i_cast_pe                 (cast_data_i_1_6),
    .ready_o_cast_pe                (cast_ready_o_1_6),
    .valid_o_cast_pe                (cast_valid_o_1_6),
    .data_o_cast_pe                 (cast_data_o_1_6),
    .ready_i_cast_pe                (cast_ready_i_1_6),

    .valid_i_merge_pe               (merge_valid_i_1_6),
    .data_i_merge_pe                (merge_data_i_1_6),
    .ready_o_merge_pe               (merge_ready_o_1_6),
    .valid_o_merge_pe               (merge_valid_o_1_6),
    .data_o_merge_pe                (merge_data_o_1_6),
    .ready_i_merge_pe               (merge_ready_i_1_6),

    .valid_i_gather_pe              (gather_valid_i_1_6),
    .data_i_gather_pe               (gather_data_i_1_6),
    .ready_o_gather_pe              (gather_ready_o_1_6),
    .valid_o_gather_pe              (gather_valid_o_1_6),
    .data_o_gather_pe               (gather_data_o_1_6),
    .ready_i_gather_pe              (gather_ready_i_1_6),

    .credit_upd                     (credit_upd[1][6])
);


network_interface #(
    .cast_out                       (cast_out_1_7),
    .gather_out                     (gather_out_1_7),
    .cast_sid                       (cast_sid_1_7),
    .gather_sid                     (gather_sid_1_7)
)ni_1_7(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[1][7]),
    .data_i_cast_nw                 (data_o_cast_nw[1][7]),
    .ready_o_cast_nw                (ready_i_cast_nw[1][7]),
    .valid_o_cast_nw                (valid_i_cast_nw[1][7]),
    .data_o_cast_nw                 (data_i_cast_nw[1][7]),
    .ready_i_cast_nw                (ready_o_cast_nw[1][7]),

    .valid_i_gather_nw              (valid_o_gather_nw[1][7]),
    .data_i_gather_nw               (data_o_gather_nw[1][7]),
    .ready_o_gather_nw              (ready_i_gather_nw[1][7]),
    .valid_o_gather_nw              (valid_i_gather_nw[1][7]),
    .data_o_gather_nw               (data_i_gather_nw[1][7]),
    .ready_i_gather_nw              (ready_o_gather_nw[1][7]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[1][7]),
    .data_i_merge_nw                (data_o_merge_nw[1][7]),
    .ready_o_merge_nw               (ready_i_merge_nw[1][7]),
    .valid_o_merge_nw               (valid_i_merge_nw[1][7]),
    .data_o_merge_nw                (data_i_merge_nw[1][7]),
    .ready_i_merge_nw               (ready_o_merge_nw[1][7]),

    .valid_i_cast_pe                (cast_valid_i_1_7),
    .data_i_cast_pe                 (cast_data_i_1_7),
    .ready_o_cast_pe                (cast_ready_o_1_7),
    .valid_o_cast_pe                (cast_valid_o_1_7),
    .data_o_cast_pe                 (cast_data_o_1_7),
    .ready_i_cast_pe                (cast_ready_i_1_7),

    .valid_i_merge_pe               (merge_valid_i_1_7),
    .data_i_merge_pe                (merge_data_i_1_7),
    .ready_o_merge_pe               (merge_ready_o_1_7),
    .valid_o_merge_pe               (merge_valid_o_1_7),
    .data_o_merge_pe                (merge_data_o_1_7),
    .ready_i_merge_pe               (merge_ready_i_1_7),

    .valid_i_gather_pe              (gather_valid_i_1_7),
    .data_i_gather_pe               (gather_data_i_1_7),
    .ready_o_gather_pe              (gather_ready_o_1_7),
    .valid_o_gather_pe              (gather_valid_o_1_7),
    .data_o_gather_pe               (gather_data_o_1_7),
    .ready_i_gather_pe              (gather_ready_i_1_7),

    .credit_upd                     (credit_upd[1][7])
);


network_interface #(
    .cast_out                       (cast_out_1_8),
    .gather_out                     (gather_out_1_8),
    .cast_sid                       (cast_sid_1_8),
    .gather_sid                     (gather_sid_1_8)
)ni_1_8(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[1][8]),
    .data_i_cast_nw                 (data_o_cast_nw[1][8]),
    .ready_o_cast_nw                (ready_i_cast_nw[1][8]),
    .valid_o_cast_nw                (valid_i_cast_nw[1][8]),
    .data_o_cast_nw                 (data_i_cast_nw[1][8]),
    .ready_i_cast_nw                (ready_o_cast_nw[1][8]),

    .valid_i_gather_nw              (valid_o_gather_nw[1][8]),
    .data_i_gather_nw               (data_o_gather_nw[1][8]),
    .ready_o_gather_nw              (ready_i_gather_nw[1][8]),
    .valid_o_gather_nw              (valid_i_gather_nw[1][8]),
    .data_o_gather_nw               (data_i_gather_nw[1][8]),
    .ready_i_gather_nw              (ready_o_gather_nw[1][8]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[1][8]),
    .data_i_merge_nw                (data_o_merge_nw[1][8]),
    .ready_o_merge_nw               (ready_i_merge_nw[1][8]),
    .valid_o_merge_nw               (valid_i_merge_nw[1][8]),
    .data_o_merge_nw                (data_i_merge_nw[1][8]),
    .ready_i_merge_nw               (ready_o_merge_nw[1][8]),

    .valid_i_cast_pe                (cast_valid_i_1_8),
    .data_i_cast_pe                 (cast_data_i_1_8),
    .ready_o_cast_pe                (cast_ready_o_1_8),
    .valid_o_cast_pe                (cast_valid_o_1_8),
    .data_o_cast_pe                 (cast_data_o_1_8),
    .ready_i_cast_pe                (cast_ready_i_1_8),

    .valid_i_merge_pe               (merge_valid_i_1_8),
    .data_i_merge_pe                (merge_data_i_1_8),
    .ready_o_merge_pe               (merge_ready_o_1_8),
    .valid_o_merge_pe               (merge_valid_o_1_8),
    .data_o_merge_pe                (merge_data_o_1_8),
    .ready_i_merge_pe               (merge_ready_i_1_8),

    .valid_i_gather_pe              (gather_valid_i_1_8),
    .data_i_gather_pe               (gather_data_i_1_8),
    .ready_o_gather_pe              (gather_ready_o_1_8),
    .valid_o_gather_pe              (gather_valid_o_1_8),
    .data_o_gather_pe               (gather_data_o_1_8),
    .ready_i_gather_pe              (gather_ready_i_1_8),

    .credit_upd                     (credit_upd[1][8])
);


network_interface #(
    .cast_out                       (cast_out_1_9),
    .gather_out                     (gather_out_1_9),
    .cast_sid                       (cast_sid_1_9),
    .gather_sid                     (gather_sid_1_9)
)ni_1_9(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[1][9]),
    .data_i_cast_nw                 (data_o_cast_nw[1][9]),
    .ready_o_cast_nw                (ready_i_cast_nw[1][9]),
    .valid_o_cast_nw                (valid_i_cast_nw[1][9]),
    .data_o_cast_nw                 (data_i_cast_nw[1][9]),
    .ready_i_cast_nw                (ready_o_cast_nw[1][9]),

    .valid_i_gather_nw              (valid_o_gather_nw[1][9]),
    .data_i_gather_nw               (data_o_gather_nw[1][9]),
    .ready_o_gather_nw              (ready_i_gather_nw[1][9]),
    .valid_o_gather_nw              (valid_i_gather_nw[1][9]),
    .data_o_gather_nw               (data_i_gather_nw[1][9]),
    .ready_i_gather_nw              (ready_o_gather_nw[1][9]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[1][9]),
    .data_i_merge_nw                (data_o_merge_nw[1][9]),
    .ready_o_merge_nw               (ready_i_merge_nw[1][9]),
    .valid_o_merge_nw               (valid_i_merge_nw[1][9]),
    .data_o_merge_nw                (data_i_merge_nw[1][9]),
    .ready_i_merge_nw               (ready_o_merge_nw[1][9]),

    .valid_i_cast_pe                (cast_valid_i_1_9),
    .data_i_cast_pe                 (cast_data_i_1_9),
    .ready_o_cast_pe                (cast_ready_o_1_9),
    .valid_o_cast_pe                (cast_valid_o_1_9),
    .data_o_cast_pe                 (cast_data_o_1_9),
    .ready_i_cast_pe                (cast_ready_i_1_9),

    .valid_i_merge_pe               (merge_valid_i_1_9),
    .data_i_merge_pe                (merge_data_i_1_9),
    .ready_o_merge_pe               (merge_ready_o_1_9),
    .valid_o_merge_pe               (merge_valid_o_1_9),
    .data_o_merge_pe                (merge_data_o_1_9),
    .ready_i_merge_pe               (merge_ready_i_1_9),

    .valid_i_gather_pe              (gather_valid_i_1_9),
    .data_i_gather_pe               (gather_data_i_1_9),
    .ready_o_gather_pe              (gather_ready_o_1_9),
    .valid_o_gather_pe              (gather_valid_o_1_9),
    .data_o_gather_pe               (gather_data_o_1_9),
    .ready_i_gather_pe              (gather_ready_i_1_9),

    .credit_upd                     (credit_upd[1][9])
);


network_interface #(
    .cast_out                       (cast_out_2_0),
    .gather_out                     (gather_out_2_0),
    .cast_sid                       (cast_sid_2_0),
    .gather_sid                     (gather_sid_2_0)
)ni_2_0(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[2][0]),
    .data_i_cast_nw                 (data_o_cast_nw[2][0]),
    .ready_o_cast_nw                (ready_i_cast_nw[2][0]),
    .valid_o_cast_nw                (valid_i_cast_nw[2][0]),
    .data_o_cast_nw                 (data_i_cast_nw[2][0]),
    .ready_i_cast_nw                (ready_o_cast_nw[2][0]),

    .valid_i_gather_nw              (valid_o_gather_nw[2][0]),
    .data_i_gather_nw               (data_o_gather_nw[2][0]),
    .ready_o_gather_nw              (ready_i_gather_nw[2][0]),
    .valid_o_gather_nw              (valid_i_gather_nw[2][0]),
    .data_o_gather_nw               (data_i_gather_nw[2][0]),
    .ready_i_gather_nw              (ready_o_gather_nw[2][0]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[2][0]),
    .data_i_merge_nw                (data_o_merge_nw[2][0]),
    .ready_o_merge_nw               (ready_i_merge_nw[2][0]),
    .valid_o_merge_nw               (valid_i_merge_nw[2][0]),
    .data_o_merge_nw                (data_i_merge_nw[2][0]),
    .ready_i_merge_nw               (ready_o_merge_nw[2][0]),

    .valid_i_cast_pe                (cast_valid_i_2_0),
    .data_i_cast_pe                 (cast_data_i_2_0),
    .ready_o_cast_pe                (cast_ready_o_2_0),
    .valid_o_cast_pe                (cast_valid_o_2_0),
    .data_o_cast_pe                 (cast_data_o_2_0),
    .ready_i_cast_pe                (cast_ready_i_2_0),

    .valid_i_merge_pe               (merge_valid_i_2_0),
    .data_i_merge_pe                (merge_data_i_2_0),
    .ready_o_merge_pe               (merge_ready_o_2_0),
    .valid_o_merge_pe               (merge_valid_o_2_0),
    .data_o_merge_pe                (merge_data_o_2_0),
    .ready_i_merge_pe               (merge_ready_i_2_0),

    .valid_i_gather_pe              (gather_valid_i_2_0),
    .data_i_gather_pe               (gather_data_i_2_0),
    .ready_o_gather_pe              (gather_ready_o_2_0),
    .valid_o_gather_pe              (gather_valid_o_2_0),
    .data_o_gather_pe               (gather_data_o_2_0),
    .ready_i_gather_pe              (gather_ready_i_2_0),

    .credit_upd                     (credit_upd[2][0])
);


network_interface #(
    .cast_out                       (cast_out_2_1),
    .gather_out                     (gather_out_2_1),
    .cast_sid                       (cast_sid_2_1),
    .gather_sid                     (gather_sid_2_1)
)ni_2_1(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[2][1]),
    .data_i_cast_nw                 (data_o_cast_nw[2][1]),
    .ready_o_cast_nw                (ready_i_cast_nw[2][1]),
    .valid_o_cast_nw                (valid_i_cast_nw[2][1]),
    .data_o_cast_nw                 (data_i_cast_nw[2][1]),
    .ready_i_cast_nw                (ready_o_cast_nw[2][1]),

    .valid_i_gather_nw              (valid_o_gather_nw[2][1]),
    .data_i_gather_nw               (data_o_gather_nw[2][1]),
    .ready_o_gather_nw              (ready_i_gather_nw[2][1]),
    .valid_o_gather_nw              (valid_i_gather_nw[2][1]),
    .data_o_gather_nw               (data_i_gather_nw[2][1]),
    .ready_i_gather_nw              (ready_o_gather_nw[2][1]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[2][1]),
    .data_i_merge_nw                (data_o_merge_nw[2][1]),
    .ready_o_merge_nw               (ready_i_merge_nw[2][1]),
    .valid_o_merge_nw               (valid_i_merge_nw[2][1]),
    .data_o_merge_nw                (data_i_merge_nw[2][1]),
    .ready_i_merge_nw               (ready_o_merge_nw[2][1]),

    .valid_i_cast_pe                (cast_valid_i_2_1),
    .data_i_cast_pe                 (cast_data_i_2_1),
    .ready_o_cast_pe                (cast_ready_o_2_1),
    .valid_o_cast_pe                (cast_valid_o_2_1),
    .data_o_cast_pe                 (cast_data_o_2_1),
    .ready_i_cast_pe                (cast_ready_i_2_1),

    .valid_i_merge_pe               (merge_valid_i_2_1),
    .data_i_merge_pe                (merge_data_i_2_1),
    .ready_o_merge_pe               (merge_ready_o_2_1),
    .valid_o_merge_pe               (merge_valid_o_2_1),
    .data_o_merge_pe                (merge_data_o_2_1),
    .ready_i_merge_pe               (merge_ready_i_2_1),

    .valid_i_gather_pe              (gather_valid_i_2_1),
    .data_i_gather_pe               (gather_data_i_2_1),
    .ready_o_gather_pe              (gather_ready_o_2_1),
    .valid_o_gather_pe              (gather_valid_o_2_1),
    .data_o_gather_pe               (gather_data_o_2_1),
    .ready_i_gather_pe              (gather_ready_i_2_1),

    .credit_upd                     (credit_upd[2][1])
);


network_interface #(
    .cast_out                       (cast_out_2_2),
    .gather_out                     (gather_out_2_2),
    .cast_sid                       (cast_sid_2_2),
    .gather_sid                     (gather_sid_2_2)
)ni_2_2(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[2][2]),
    .data_i_cast_nw                 (data_o_cast_nw[2][2]),
    .ready_o_cast_nw                (ready_i_cast_nw[2][2]),
    .valid_o_cast_nw                (valid_i_cast_nw[2][2]),
    .data_o_cast_nw                 (data_i_cast_nw[2][2]),
    .ready_i_cast_nw                (ready_o_cast_nw[2][2]),

    .valid_i_gather_nw              (valid_o_gather_nw[2][2]),
    .data_i_gather_nw               (data_o_gather_nw[2][2]),
    .ready_o_gather_nw              (ready_i_gather_nw[2][2]),
    .valid_o_gather_nw              (valid_i_gather_nw[2][2]),
    .data_o_gather_nw               (data_i_gather_nw[2][2]),
    .ready_i_gather_nw              (ready_o_gather_nw[2][2]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[2][2]),
    .data_i_merge_nw                (data_o_merge_nw[2][2]),
    .ready_o_merge_nw               (ready_i_merge_nw[2][2]),
    .valid_o_merge_nw               (valid_i_merge_nw[2][2]),
    .data_o_merge_nw                (data_i_merge_nw[2][2]),
    .ready_i_merge_nw               (ready_o_merge_nw[2][2]),

    .valid_i_cast_pe                (cast_valid_i_2_2),
    .data_i_cast_pe                 (cast_data_i_2_2),
    .ready_o_cast_pe                (cast_ready_o_2_2),
    .valid_o_cast_pe                (cast_valid_o_2_2),
    .data_o_cast_pe                 (cast_data_o_2_2),
    .ready_i_cast_pe                (cast_ready_i_2_2),

    .valid_i_merge_pe               (merge_valid_i_2_2),
    .data_i_merge_pe                (merge_data_i_2_2),
    .ready_o_merge_pe               (merge_ready_o_2_2),
    .valid_o_merge_pe               (merge_valid_o_2_2),
    .data_o_merge_pe                (merge_data_o_2_2),
    .ready_i_merge_pe               (merge_ready_i_2_2),

    .valid_i_gather_pe              (gather_valid_i_2_2),
    .data_i_gather_pe               (gather_data_i_2_2),
    .ready_o_gather_pe              (gather_ready_o_2_2),
    .valid_o_gather_pe              (gather_valid_o_2_2),
    .data_o_gather_pe               (gather_data_o_2_2),
    .ready_i_gather_pe              (gather_ready_i_2_2),

    .credit_upd                     (credit_upd[2][2])
);


network_interface #(
    .cast_out                       (cast_out_2_3),
    .gather_out                     (gather_out_2_3),
    .cast_sid                       (cast_sid_2_3),
    .gather_sid                     (gather_sid_2_3)
)ni_2_3(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[2][3]),
    .data_i_cast_nw                 (data_o_cast_nw[2][3]),
    .ready_o_cast_nw                (ready_i_cast_nw[2][3]),
    .valid_o_cast_nw                (valid_i_cast_nw[2][3]),
    .data_o_cast_nw                 (data_i_cast_nw[2][3]),
    .ready_i_cast_nw                (ready_o_cast_nw[2][3]),

    .valid_i_gather_nw              (valid_o_gather_nw[2][3]),
    .data_i_gather_nw               (data_o_gather_nw[2][3]),
    .ready_o_gather_nw              (ready_i_gather_nw[2][3]),
    .valid_o_gather_nw              (valid_i_gather_nw[2][3]),
    .data_o_gather_nw               (data_i_gather_nw[2][3]),
    .ready_i_gather_nw              (ready_o_gather_nw[2][3]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[2][3]),
    .data_i_merge_nw                (data_o_merge_nw[2][3]),
    .ready_o_merge_nw               (ready_i_merge_nw[2][3]),
    .valid_o_merge_nw               (valid_i_merge_nw[2][3]),
    .data_o_merge_nw                (data_i_merge_nw[2][3]),
    .ready_i_merge_nw               (ready_o_merge_nw[2][3]),

    .valid_i_cast_pe                (cast_valid_i_2_3),
    .data_i_cast_pe                 (cast_data_i_2_3),
    .ready_o_cast_pe                (cast_ready_o_2_3),
    .valid_o_cast_pe                (cast_valid_o_2_3),
    .data_o_cast_pe                 (cast_data_o_2_3),
    .ready_i_cast_pe                (cast_ready_i_2_3),

    .valid_i_merge_pe               (merge_valid_i_2_3),
    .data_i_merge_pe                (merge_data_i_2_3),
    .ready_o_merge_pe               (merge_ready_o_2_3),
    .valid_o_merge_pe               (merge_valid_o_2_3),
    .data_o_merge_pe                (merge_data_o_2_3),
    .ready_i_merge_pe               (merge_ready_i_2_3),

    .valid_i_gather_pe              (gather_valid_i_2_3),
    .data_i_gather_pe               (gather_data_i_2_3),
    .ready_o_gather_pe              (gather_ready_o_2_3),
    .valid_o_gather_pe              (gather_valid_o_2_3),
    .data_o_gather_pe               (gather_data_o_2_3),
    .ready_i_gather_pe              (gather_ready_i_2_3),

    .credit_upd                     (credit_upd[2][3])
);


network_interface #(
    .cast_out                       (cast_out_2_4),
    .gather_out                     (gather_out_2_4),
    .cast_sid                       (cast_sid_2_4),
    .gather_sid                     (gather_sid_2_4)
)ni_2_4(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[2][4]),
    .data_i_cast_nw                 (data_o_cast_nw[2][4]),
    .ready_o_cast_nw                (ready_i_cast_nw[2][4]),
    .valid_o_cast_nw                (valid_i_cast_nw[2][4]),
    .data_o_cast_nw                 (data_i_cast_nw[2][4]),
    .ready_i_cast_nw                (ready_o_cast_nw[2][4]),

    .valid_i_gather_nw              (valid_o_gather_nw[2][4]),
    .data_i_gather_nw               (data_o_gather_nw[2][4]),
    .ready_o_gather_nw              (ready_i_gather_nw[2][4]),
    .valid_o_gather_nw              (valid_i_gather_nw[2][4]),
    .data_o_gather_nw               (data_i_gather_nw[2][4]),
    .ready_i_gather_nw              (ready_o_gather_nw[2][4]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[2][4]),
    .data_i_merge_nw                (data_o_merge_nw[2][4]),
    .ready_o_merge_nw               (ready_i_merge_nw[2][4]),
    .valid_o_merge_nw               (valid_i_merge_nw[2][4]),
    .data_o_merge_nw                (data_i_merge_nw[2][4]),
    .ready_i_merge_nw               (ready_o_merge_nw[2][4]),

    .valid_i_cast_pe                (cast_valid_i_2_4),
    .data_i_cast_pe                 (cast_data_i_2_4),
    .ready_o_cast_pe                (cast_ready_o_2_4),
    .valid_o_cast_pe                (cast_valid_o_2_4),
    .data_o_cast_pe                 (cast_data_o_2_4),
    .ready_i_cast_pe                (cast_ready_i_2_4),

    .valid_i_merge_pe               (merge_valid_i_2_4),
    .data_i_merge_pe                (merge_data_i_2_4),
    .ready_o_merge_pe               (merge_ready_o_2_4),
    .valid_o_merge_pe               (merge_valid_o_2_4),
    .data_o_merge_pe                (merge_data_o_2_4),
    .ready_i_merge_pe               (merge_ready_i_2_4),

    .valid_i_gather_pe              (gather_valid_i_2_4),
    .data_i_gather_pe               (gather_data_i_2_4),
    .ready_o_gather_pe              (gather_ready_o_2_4),
    .valid_o_gather_pe              (gather_valid_o_2_4),
    .data_o_gather_pe               (gather_data_o_2_4),
    .ready_i_gather_pe              (gather_ready_i_2_4),

    .credit_upd                     (credit_upd[2][4])
);


network_interface #(
    .cast_out                       (cast_out_2_5),
    .gather_out                     (gather_out_2_5),
    .cast_sid                       (cast_sid_2_5),
    .gather_sid                     (gather_sid_2_5)
)ni_2_5(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[2][5]),
    .data_i_cast_nw                 (data_o_cast_nw[2][5]),
    .ready_o_cast_nw                (ready_i_cast_nw[2][5]),
    .valid_o_cast_nw                (valid_i_cast_nw[2][5]),
    .data_o_cast_nw                 (data_i_cast_nw[2][5]),
    .ready_i_cast_nw                (ready_o_cast_nw[2][5]),

    .valid_i_gather_nw              (valid_o_gather_nw[2][5]),
    .data_i_gather_nw               (data_o_gather_nw[2][5]),
    .ready_o_gather_nw              (ready_i_gather_nw[2][5]),
    .valid_o_gather_nw              (valid_i_gather_nw[2][5]),
    .data_o_gather_nw               (data_i_gather_nw[2][5]),
    .ready_i_gather_nw              (ready_o_gather_nw[2][5]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[2][5]),
    .data_i_merge_nw                (data_o_merge_nw[2][5]),
    .ready_o_merge_nw               (ready_i_merge_nw[2][5]),
    .valid_o_merge_nw               (valid_i_merge_nw[2][5]),
    .data_o_merge_nw                (data_i_merge_nw[2][5]),
    .ready_i_merge_nw               (ready_o_merge_nw[2][5]),

    .valid_i_cast_pe                (cast_valid_i_2_5),
    .data_i_cast_pe                 (cast_data_i_2_5),
    .ready_o_cast_pe                (cast_ready_o_2_5),
    .valid_o_cast_pe                (cast_valid_o_2_5),
    .data_o_cast_pe                 (cast_data_o_2_5),
    .ready_i_cast_pe                (cast_ready_i_2_5),

    .valid_i_merge_pe               (merge_valid_i_2_5),
    .data_i_merge_pe                (merge_data_i_2_5),
    .ready_o_merge_pe               (merge_ready_o_2_5),
    .valid_o_merge_pe               (merge_valid_o_2_5),
    .data_o_merge_pe                (merge_data_o_2_5),
    .ready_i_merge_pe               (merge_ready_i_2_5),

    .valid_i_gather_pe              (gather_valid_i_2_5),
    .data_i_gather_pe               (gather_data_i_2_5),
    .ready_o_gather_pe              (gather_ready_o_2_5),
    .valid_o_gather_pe              (gather_valid_o_2_5),
    .data_o_gather_pe               (gather_data_o_2_5),
    .ready_i_gather_pe              (gather_ready_i_2_5),

    .credit_upd                     (credit_upd[2][5])
);


network_interface #(
    .cast_out                       (cast_out_2_6),
    .gather_out                     (gather_out_2_6),
    .cast_sid                       (cast_sid_2_6),
    .gather_sid                     (gather_sid_2_6)
)ni_2_6(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[2][6]),
    .data_i_cast_nw                 (data_o_cast_nw[2][6]),
    .ready_o_cast_nw                (ready_i_cast_nw[2][6]),
    .valid_o_cast_nw                (valid_i_cast_nw[2][6]),
    .data_o_cast_nw                 (data_i_cast_nw[2][6]),
    .ready_i_cast_nw                (ready_o_cast_nw[2][6]),

    .valid_i_gather_nw              (valid_o_gather_nw[2][6]),
    .data_i_gather_nw               (data_o_gather_nw[2][6]),
    .ready_o_gather_nw              (ready_i_gather_nw[2][6]),
    .valid_o_gather_nw              (valid_i_gather_nw[2][6]),
    .data_o_gather_nw               (data_i_gather_nw[2][6]),
    .ready_i_gather_nw              (ready_o_gather_nw[2][6]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[2][6]),
    .data_i_merge_nw                (data_o_merge_nw[2][6]),
    .ready_o_merge_nw               (ready_i_merge_nw[2][6]),
    .valid_o_merge_nw               (valid_i_merge_nw[2][6]),
    .data_o_merge_nw                (data_i_merge_nw[2][6]),
    .ready_i_merge_nw               (ready_o_merge_nw[2][6]),

    .valid_i_cast_pe                (cast_valid_i_2_6),
    .data_i_cast_pe                 (cast_data_i_2_6),
    .ready_o_cast_pe                (cast_ready_o_2_6),
    .valid_o_cast_pe                (cast_valid_o_2_6),
    .data_o_cast_pe                 (cast_data_o_2_6),
    .ready_i_cast_pe                (cast_ready_i_2_6),

    .valid_i_merge_pe               (merge_valid_i_2_6),
    .data_i_merge_pe                (merge_data_i_2_6),
    .ready_o_merge_pe               (merge_ready_o_2_6),
    .valid_o_merge_pe               (merge_valid_o_2_6),
    .data_o_merge_pe                (merge_data_o_2_6),
    .ready_i_merge_pe               (merge_ready_i_2_6),

    .valid_i_gather_pe              (gather_valid_i_2_6),
    .data_i_gather_pe               (gather_data_i_2_6),
    .ready_o_gather_pe              (gather_ready_o_2_6),
    .valid_o_gather_pe              (gather_valid_o_2_6),
    .data_o_gather_pe               (gather_data_o_2_6),
    .ready_i_gather_pe              (gather_ready_i_2_6),

    .credit_upd                     (credit_upd[2][6])
);


network_interface #(
    .cast_out                       (cast_out_2_7),
    .gather_out                     (gather_out_2_7),
    .cast_sid                       (cast_sid_2_7),
    .gather_sid                     (gather_sid_2_7)
)ni_2_7(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[2][7]),
    .data_i_cast_nw                 (data_o_cast_nw[2][7]),
    .ready_o_cast_nw                (ready_i_cast_nw[2][7]),
    .valid_o_cast_nw                (valid_i_cast_nw[2][7]),
    .data_o_cast_nw                 (data_i_cast_nw[2][7]),
    .ready_i_cast_nw                (ready_o_cast_nw[2][7]),

    .valid_i_gather_nw              (valid_o_gather_nw[2][7]),
    .data_i_gather_nw               (data_o_gather_nw[2][7]),
    .ready_o_gather_nw              (ready_i_gather_nw[2][7]),
    .valid_o_gather_nw              (valid_i_gather_nw[2][7]),
    .data_o_gather_nw               (data_i_gather_nw[2][7]),
    .ready_i_gather_nw              (ready_o_gather_nw[2][7]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[2][7]),
    .data_i_merge_nw                (data_o_merge_nw[2][7]),
    .ready_o_merge_nw               (ready_i_merge_nw[2][7]),
    .valid_o_merge_nw               (valid_i_merge_nw[2][7]),
    .data_o_merge_nw                (data_i_merge_nw[2][7]),
    .ready_i_merge_nw               (ready_o_merge_nw[2][7]),

    .valid_i_cast_pe                (cast_valid_i_2_7),
    .data_i_cast_pe                 (cast_data_i_2_7),
    .ready_o_cast_pe                (cast_ready_o_2_7),
    .valid_o_cast_pe                (cast_valid_o_2_7),
    .data_o_cast_pe                 (cast_data_o_2_7),
    .ready_i_cast_pe                (cast_ready_i_2_7),

    .valid_i_merge_pe               (merge_valid_i_2_7),
    .data_i_merge_pe                (merge_data_i_2_7),
    .ready_o_merge_pe               (merge_ready_o_2_7),
    .valid_o_merge_pe               (merge_valid_o_2_7),
    .data_o_merge_pe                (merge_data_o_2_7),
    .ready_i_merge_pe               (merge_ready_i_2_7),

    .valid_i_gather_pe              (gather_valid_i_2_7),
    .data_i_gather_pe               (gather_data_i_2_7),
    .ready_o_gather_pe              (gather_ready_o_2_7),
    .valid_o_gather_pe              (gather_valid_o_2_7),
    .data_o_gather_pe               (gather_data_o_2_7),
    .ready_i_gather_pe              (gather_ready_i_2_7),

    .credit_upd                     (credit_upd[2][7])
);


network_interface #(
    .cast_out                       (cast_out_2_8),
    .gather_out                     (gather_out_2_8),
    .cast_sid                       (cast_sid_2_8),
    .gather_sid                     (gather_sid_2_8)
)ni_2_8(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[2][8]),
    .data_i_cast_nw                 (data_o_cast_nw[2][8]),
    .ready_o_cast_nw                (ready_i_cast_nw[2][8]),
    .valid_o_cast_nw                (valid_i_cast_nw[2][8]),
    .data_o_cast_nw                 (data_i_cast_nw[2][8]),
    .ready_i_cast_nw                (ready_o_cast_nw[2][8]),

    .valid_i_gather_nw              (valid_o_gather_nw[2][8]),
    .data_i_gather_nw               (data_o_gather_nw[2][8]),
    .ready_o_gather_nw              (ready_i_gather_nw[2][8]),
    .valid_o_gather_nw              (valid_i_gather_nw[2][8]),
    .data_o_gather_nw               (data_i_gather_nw[2][8]),
    .ready_i_gather_nw              (ready_o_gather_nw[2][8]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[2][8]),
    .data_i_merge_nw                (data_o_merge_nw[2][8]),
    .ready_o_merge_nw               (ready_i_merge_nw[2][8]),
    .valid_o_merge_nw               (valid_i_merge_nw[2][8]),
    .data_o_merge_nw                (data_i_merge_nw[2][8]),
    .ready_i_merge_nw               (ready_o_merge_nw[2][8]),

    .valid_i_cast_pe                (cast_valid_i_2_8),
    .data_i_cast_pe                 (cast_data_i_2_8),
    .ready_o_cast_pe                (cast_ready_o_2_8),
    .valid_o_cast_pe                (cast_valid_o_2_8),
    .data_o_cast_pe                 (cast_data_o_2_8),
    .ready_i_cast_pe                (cast_ready_i_2_8),

    .valid_i_merge_pe               (merge_valid_i_2_8),
    .data_i_merge_pe                (merge_data_i_2_8),
    .ready_o_merge_pe               (merge_ready_o_2_8),
    .valid_o_merge_pe               (merge_valid_o_2_8),
    .data_o_merge_pe                (merge_data_o_2_8),
    .ready_i_merge_pe               (merge_ready_i_2_8),

    .valid_i_gather_pe              (gather_valid_i_2_8),
    .data_i_gather_pe               (gather_data_i_2_8),
    .ready_o_gather_pe              (gather_ready_o_2_8),
    .valid_o_gather_pe              (gather_valid_o_2_8),
    .data_o_gather_pe               (gather_data_o_2_8),
    .ready_i_gather_pe              (gather_ready_i_2_8),

    .credit_upd                     (credit_upd[2][8])
);


network_interface #(
    .cast_out                       (cast_out_2_9),
    .gather_out                     (gather_out_2_9),
    .cast_sid                       (cast_sid_2_9),
    .gather_sid                     (gather_sid_2_9)
)ni_2_9(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[2][9]),
    .data_i_cast_nw                 (data_o_cast_nw[2][9]),
    .ready_o_cast_nw                (ready_i_cast_nw[2][9]),
    .valid_o_cast_nw                (valid_i_cast_nw[2][9]),
    .data_o_cast_nw                 (data_i_cast_nw[2][9]),
    .ready_i_cast_nw                (ready_o_cast_nw[2][9]),

    .valid_i_gather_nw              (valid_o_gather_nw[2][9]),
    .data_i_gather_nw               (data_o_gather_nw[2][9]),
    .ready_o_gather_nw              (ready_i_gather_nw[2][9]),
    .valid_o_gather_nw              (valid_i_gather_nw[2][9]),
    .data_o_gather_nw               (data_i_gather_nw[2][9]),
    .ready_i_gather_nw              (ready_o_gather_nw[2][9]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[2][9]),
    .data_i_merge_nw                (data_o_merge_nw[2][9]),
    .ready_o_merge_nw               (ready_i_merge_nw[2][9]),
    .valid_o_merge_nw               (valid_i_merge_nw[2][9]),
    .data_o_merge_nw                (data_i_merge_nw[2][9]),
    .ready_i_merge_nw               (ready_o_merge_nw[2][9]),

    .valid_i_cast_pe                (cast_valid_i_2_9),
    .data_i_cast_pe                 (cast_data_i_2_9),
    .ready_o_cast_pe                (cast_ready_o_2_9),
    .valid_o_cast_pe                (cast_valid_o_2_9),
    .data_o_cast_pe                 (cast_data_o_2_9),
    .ready_i_cast_pe                (cast_ready_i_2_9),

    .valid_i_merge_pe               (merge_valid_i_2_9),
    .data_i_merge_pe                (merge_data_i_2_9),
    .ready_o_merge_pe               (merge_ready_o_2_9),
    .valid_o_merge_pe               (merge_valid_o_2_9),
    .data_o_merge_pe                (merge_data_o_2_9),
    .ready_i_merge_pe               (merge_ready_i_2_9),

    .valid_i_gather_pe              (gather_valid_i_2_9),
    .data_i_gather_pe               (gather_data_i_2_9),
    .ready_o_gather_pe              (gather_ready_o_2_9),
    .valid_o_gather_pe              (gather_valid_o_2_9),
    .data_o_gather_pe               (gather_data_o_2_9),
    .ready_i_gather_pe              (gather_ready_i_2_9),

    .credit_upd                     (credit_upd[2][9])
);


network_interface #(
    .cast_out                       (cast_out_3_0),
    .gather_out                     (gather_out_3_0),
    .cast_sid                       (cast_sid_3_0),
    .gather_sid                     (gather_sid_3_0)
)ni_3_0(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[3][0]),
    .data_i_cast_nw                 (data_o_cast_nw[3][0]),
    .ready_o_cast_nw                (ready_i_cast_nw[3][0]),
    .valid_o_cast_nw                (valid_i_cast_nw[3][0]),
    .data_o_cast_nw                 (data_i_cast_nw[3][0]),
    .ready_i_cast_nw                (ready_o_cast_nw[3][0]),

    .valid_i_gather_nw              (valid_o_gather_nw[3][0]),
    .data_i_gather_nw               (data_o_gather_nw[3][0]),
    .ready_o_gather_nw              (ready_i_gather_nw[3][0]),
    .valid_o_gather_nw              (valid_i_gather_nw[3][0]),
    .data_o_gather_nw               (data_i_gather_nw[3][0]),
    .ready_i_gather_nw              (ready_o_gather_nw[3][0]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[3][0]),
    .data_i_merge_nw                (data_o_merge_nw[3][0]),
    .ready_o_merge_nw               (ready_i_merge_nw[3][0]),
    .valid_o_merge_nw               (valid_i_merge_nw[3][0]),
    .data_o_merge_nw                (data_i_merge_nw[3][0]),
    .ready_i_merge_nw               (ready_o_merge_nw[3][0]),

    .valid_i_cast_pe                (cast_valid_i_3_0),
    .data_i_cast_pe                 (cast_data_i_3_0),
    .ready_o_cast_pe                (cast_ready_o_3_0),
    .valid_o_cast_pe                (cast_valid_o_3_0),
    .data_o_cast_pe                 (cast_data_o_3_0),
    .ready_i_cast_pe                (cast_ready_i_3_0),

    .valid_i_merge_pe               (merge_valid_i_3_0),
    .data_i_merge_pe                (merge_data_i_3_0),
    .ready_o_merge_pe               (merge_ready_o_3_0),
    .valid_o_merge_pe               (merge_valid_o_3_0),
    .data_o_merge_pe                (merge_data_o_3_0),
    .ready_i_merge_pe               (merge_ready_i_3_0),

    .valid_i_gather_pe              (gather_valid_i_3_0),
    .data_i_gather_pe               (gather_data_i_3_0),
    .ready_o_gather_pe              (gather_ready_o_3_0),
    .valid_o_gather_pe              (gather_valid_o_3_0),
    .data_o_gather_pe               (gather_data_o_3_0),
    .ready_i_gather_pe              (gather_ready_i_3_0),

    .credit_upd                     (credit_upd[3][0])
);


network_interface #(
    .cast_out                       (cast_out_3_1),
    .gather_out                     (gather_out_3_1),
    .cast_sid                       (cast_sid_3_1),
    .gather_sid                     (gather_sid_3_1)
)ni_3_1(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[3][1]),
    .data_i_cast_nw                 (data_o_cast_nw[3][1]),
    .ready_o_cast_nw                (ready_i_cast_nw[3][1]),
    .valid_o_cast_nw                (valid_i_cast_nw[3][1]),
    .data_o_cast_nw                 (data_i_cast_nw[3][1]),
    .ready_i_cast_nw                (ready_o_cast_nw[3][1]),

    .valid_i_gather_nw              (valid_o_gather_nw[3][1]),
    .data_i_gather_nw               (data_o_gather_nw[3][1]),
    .ready_o_gather_nw              (ready_i_gather_nw[3][1]),
    .valid_o_gather_nw              (valid_i_gather_nw[3][1]),
    .data_o_gather_nw               (data_i_gather_nw[3][1]),
    .ready_i_gather_nw              (ready_o_gather_nw[3][1]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[3][1]),
    .data_i_merge_nw                (data_o_merge_nw[3][1]),
    .ready_o_merge_nw               (ready_i_merge_nw[3][1]),
    .valid_o_merge_nw               (valid_i_merge_nw[3][1]),
    .data_o_merge_nw                (data_i_merge_nw[3][1]),
    .ready_i_merge_nw               (ready_o_merge_nw[3][1]),

    .valid_i_cast_pe                (cast_valid_i_3_1),
    .data_i_cast_pe                 (cast_data_i_3_1),
    .ready_o_cast_pe                (cast_ready_o_3_1),
    .valid_o_cast_pe                (cast_valid_o_3_1),
    .data_o_cast_pe                 (cast_data_o_3_1),
    .ready_i_cast_pe                (cast_ready_i_3_1),

    .valid_i_merge_pe               (merge_valid_i_3_1),
    .data_i_merge_pe                (merge_data_i_3_1),
    .ready_o_merge_pe               (merge_ready_o_3_1),
    .valid_o_merge_pe               (merge_valid_o_3_1),
    .data_o_merge_pe                (merge_data_o_3_1),
    .ready_i_merge_pe               (merge_ready_i_3_1),

    .valid_i_gather_pe              (gather_valid_i_3_1),
    .data_i_gather_pe               (gather_data_i_3_1),
    .ready_o_gather_pe              (gather_ready_o_3_1),
    .valid_o_gather_pe              (gather_valid_o_3_1),
    .data_o_gather_pe               (gather_data_o_3_1),
    .ready_i_gather_pe              (gather_ready_i_3_1),

    .credit_upd                     (credit_upd[3][1])
);


network_interface #(
    .cast_out                       (cast_out_3_2),
    .gather_out                     (gather_out_3_2),
    .cast_sid                       (cast_sid_3_2),
    .gather_sid                     (gather_sid_3_2)
)ni_3_2(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[3][2]),
    .data_i_cast_nw                 (data_o_cast_nw[3][2]),
    .ready_o_cast_nw                (ready_i_cast_nw[3][2]),
    .valid_o_cast_nw                (valid_i_cast_nw[3][2]),
    .data_o_cast_nw                 (data_i_cast_nw[3][2]),
    .ready_i_cast_nw                (ready_o_cast_nw[3][2]),

    .valid_i_gather_nw              (valid_o_gather_nw[3][2]),
    .data_i_gather_nw               (data_o_gather_nw[3][2]),
    .ready_o_gather_nw              (ready_i_gather_nw[3][2]),
    .valid_o_gather_nw              (valid_i_gather_nw[3][2]),
    .data_o_gather_nw               (data_i_gather_nw[3][2]),
    .ready_i_gather_nw              (ready_o_gather_nw[3][2]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[3][2]),
    .data_i_merge_nw                (data_o_merge_nw[3][2]),
    .ready_o_merge_nw               (ready_i_merge_nw[3][2]),
    .valid_o_merge_nw               (valid_i_merge_nw[3][2]),
    .data_o_merge_nw                (data_i_merge_nw[3][2]),
    .ready_i_merge_nw               (ready_o_merge_nw[3][2]),

    .valid_i_cast_pe                (cast_valid_i_3_2),
    .data_i_cast_pe                 (cast_data_i_3_2),
    .ready_o_cast_pe                (cast_ready_o_3_2),
    .valid_o_cast_pe                (cast_valid_o_3_2),
    .data_o_cast_pe                 (cast_data_o_3_2),
    .ready_i_cast_pe                (cast_ready_i_3_2),

    .valid_i_merge_pe               (merge_valid_i_3_2),
    .data_i_merge_pe                (merge_data_i_3_2),
    .ready_o_merge_pe               (merge_ready_o_3_2),
    .valid_o_merge_pe               (merge_valid_o_3_2),
    .data_o_merge_pe                (merge_data_o_3_2),
    .ready_i_merge_pe               (merge_ready_i_3_2),

    .valid_i_gather_pe              (gather_valid_i_3_2),
    .data_i_gather_pe               (gather_data_i_3_2),
    .ready_o_gather_pe              (gather_ready_o_3_2),
    .valid_o_gather_pe              (gather_valid_o_3_2),
    .data_o_gather_pe               (gather_data_o_3_2),
    .ready_i_gather_pe              (gather_ready_i_3_2),

    .credit_upd                     (credit_upd[3][2])
);


network_interface #(
    .cast_out                       (cast_out_3_3),
    .gather_out                     (gather_out_3_3),
    .cast_sid                       (cast_sid_3_3),
    .gather_sid                     (gather_sid_3_3)
)ni_3_3(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[3][3]),
    .data_i_cast_nw                 (data_o_cast_nw[3][3]),
    .ready_o_cast_nw                (ready_i_cast_nw[3][3]),
    .valid_o_cast_nw                (valid_i_cast_nw[3][3]),
    .data_o_cast_nw                 (data_i_cast_nw[3][3]),
    .ready_i_cast_nw                (ready_o_cast_nw[3][3]),

    .valid_i_gather_nw              (valid_o_gather_nw[3][3]),
    .data_i_gather_nw               (data_o_gather_nw[3][3]),
    .ready_o_gather_nw              (ready_i_gather_nw[3][3]),
    .valid_o_gather_nw              (valid_i_gather_nw[3][3]),
    .data_o_gather_nw               (data_i_gather_nw[3][3]),
    .ready_i_gather_nw              (ready_o_gather_nw[3][3]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[3][3]),
    .data_i_merge_nw                (data_o_merge_nw[3][3]),
    .ready_o_merge_nw               (ready_i_merge_nw[3][3]),
    .valid_o_merge_nw               (valid_i_merge_nw[3][3]),
    .data_o_merge_nw                (data_i_merge_nw[3][3]),
    .ready_i_merge_nw               (ready_o_merge_nw[3][3]),

    .valid_i_cast_pe                (cast_valid_i_3_3),
    .data_i_cast_pe                 (cast_data_i_3_3),
    .ready_o_cast_pe                (cast_ready_o_3_3),
    .valid_o_cast_pe                (cast_valid_o_3_3),
    .data_o_cast_pe                 (cast_data_o_3_3),
    .ready_i_cast_pe                (cast_ready_i_3_3),

    .valid_i_merge_pe               (merge_valid_i_3_3),
    .data_i_merge_pe                (merge_data_i_3_3),
    .ready_o_merge_pe               (merge_ready_o_3_3),
    .valid_o_merge_pe               (merge_valid_o_3_3),
    .data_o_merge_pe                (merge_data_o_3_3),
    .ready_i_merge_pe               (merge_ready_i_3_3),

    .valid_i_gather_pe              (gather_valid_i_3_3),
    .data_i_gather_pe               (gather_data_i_3_3),
    .ready_o_gather_pe              (gather_ready_o_3_3),
    .valid_o_gather_pe              (gather_valid_o_3_3),
    .data_o_gather_pe               (gather_data_o_3_3),
    .ready_i_gather_pe              (gather_ready_i_3_3),

    .credit_upd                     (credit_upd[3][3])
);


network_interface #(
    .cast_out                       (cast_out_3_4),
    .gather_out                     (gather_out_3_4),
    .cast_sid                       (cast_sid_3_4),
    .gather_sid                     (gather_sid_3_4)
)ni_3_4(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[3][4]),
    .data_i_cast_nw                 (data_o_cast_nw[3][4]),
    .ready_o_cast_nw                (ready_i_cast_nw[3][4]),
    .valid_o_cast_nw                (valid_i_cast_nw[3][4]),
    .data_o_cast_nw                 (data_i_cast_nw[3][4]),
    .ready_i_cast_nw                (ready_o_cast_nw[3][4]),

    .valid_i_gather_nw              (valid_o_gather_nw[3][4]),
    .data_i_gather_nw               (data_o_gather_nw[3][4]),
    .ready_o_gather_nw              (ready_i_gather_nw[3][4]),
    .valid_o_gather_nw              (valid_i_gather_nw[3][4]),
    .data_o_gather_nw               (data_i_gather_nw[3][4]),
    .ready_i_gather_nw              (ready_o_gather_nw[3][4]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[3][4]),
    .data_i_merge_nw                (data_o_merge_nw[3][4]),
    .ready_o_merge_nw               (ready_i_merge_nw[3][4]),
    .valid_o_merge_nw               (valid_i_merge_nw[3][4]),
    .data_o_merge_nw                (data_i_merge_nw[3][4]),
    .ready_i_merge_nw               (ready_o_merge_nw[3][4]),

    .valid_i_cast_pe                (cast_valid_i_3_4),
    .data_i_cast_pe                 (cast_data_i_3_4),
    .ready_o_cast_pe                (cast_ready_o_3_4),
    .valid_o_cast_pe                (cast_valid_o_3_4),
    .data_o_cast_pe                 (cast_data_o_3_4),
    .ready_i_cast_pe                (cast_ready_i_3_4),

    .valid_i_merge_pe               (merge_valid_i_3_4),
    .data_i_merge_pe                (merge_data_i_3_4),
    .ready_o_merge_pe               (merge_ready_o_3_4),
    .valid_o_merge_pe               (merge_valid_o_3_4),
    .data_o_merge_pe                (merge_data_o_3_4),
    .ready_i_merge_pe               (merge_ready_i_3_4),

    .valid_i_gather_pe              (gather_valid_i_3_4),
    .data_i_gather_pe               (gather_data_i_3_4),
    .ready_o_gather_pe              (gather_ready_o_3_4),
    .valid_o_gather_pe              (gather_valid_o_3_4),
    .data_o_gather_pe               (gather_data_o_3_4),
    .ready_i_gather_pe              (gather_ready_i_3_4),

    .credit_upd                     (credit_upd[3][4])
);


network_interface #(
    .cast_out                       (cast_out_3_5),
    .gather_out                     (gather_out_3_5),
    .cast_sid                       (cast_sid_3_5),
    .gather_sid                     (gather_sid_3_5)
)ni_3_5(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[3][5]),
    .data_i_cast_nw                 (data_o_cast_nw[3][5]),
    .ready_o_cast_nw                (ready_i_cast_nw[3][5]),
    .valid_o_cast_nw                (valid_i_cast_nw[3][5]),
    .data_o_cast_nw                 (data_i_cast_nw[3][5]),
    .ready_i_cast_nw                (ready_o_cast_nw[3][5]),

    .valid_i_gather_nw              (valid_o_gather_nw[3][5]),
    .data_i_gather_nw               (data_o_gather_nw[3][5]),
    .ready_o_gather_nw              (ready_i_gather_nw[3][5]),
    .valid_o_gather_nw              (valid_i_gather_nw[3][5]),
    .data_o_gather_nw               (data_i_gather_nw[3][5]),
    .ready_i_gather_nw              (ready_o_gather_nw[3][5]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[3][5]),
    .data_i_merge_nw                (data_o_merge_nw[3][5]),
    .ready_o_merge_nw               (ready_i_merge_nw[3][5]),
    .valid_o_merge_nw               (valid_i_merge_nw[3][5]),
    .data_o_merge_nw                (data_i_merge_nw[3][5]),
    .ready_i_merge_nw               (ready_o_merge_nw[3][5]),

    .valid_i_cast_pe                (cast_valid_i_3_5),
    .data_i_cast_pe                 (cast_data_i_3_5),
    .ready_o_cast_pe                (cast_ready_o_3_5),
    .valid_o_cast_pe                (cast_valid_o_3_5),
    .data_o_cast_pe                 (cast_data_o_3_5),
    .ready_i_cast_pe                (cast_ready_i_3_5),

    .valid_i_merge_pe               (merge_valid_i_3_5),
    .data_i_merge_pe                (merge_data_i_3_5),
    .ready_o_merge_pe               (merge_ready_o_3_5),
    .valid_o_merge_pe               (merge_valid_o_3_5),
    .data_o_merge_pe                (merge_data_o_3_5),
    .ready_i_merge_pe               (merge_ready_i_3_5),

    .valid_i_gather_pe              (gather_valid_i_3_5),
    .data_i_gather_pe               (gather_data_i_3_5),
    .ready_o_gather_pe              (gather_ready_o_3_5),
    .valid_o_gather_pe              (gather_valid_o_3_5),
    .data_o_gather_pe               (gather_data_o_3_5),
    .ready_i_gather_pe              (gather_ready_i_3_5),

    .credit_upd                     (credit_upd[3][5])
);


network_interface #(
    .cast_out                       (cast_out_3_6),
    .gather_out                     (gather_out_3_6),
    .cast_sid                       (cast_sid_3_6),
    .gather_sid                     (gather_sid_3_6)
)ni_3_6(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[3][6]),
    .data_i_cast_nw                 (data_o_cast_nw[3][6]),
    .ready_o_cast_nw                (ready_i_cast_nw[3][6]),
    .valid_o_cast_nw                (valid_i_cast_nw[3][6]),
    .data_o_cast_nw                 (data_i_cast_nw[3][6]),
    .ready_i_cast_nw                (ready_o_cast_nw[3][6]),

    .valid_i_gather_nw              (valid_o_gather_nw[3][6]),
    .data_i_gather_nw               (data_o_gather_nw[3][6]),
    .ready_o_gather_nw              (ready_i_gather_nw[3][6]),
    .valid_o_gather_nw              (valid_i_gather_nw[3][6]),
    .data_o_gather_nw               (data_i_gather_nw[3][6]),
    .ready_i_gather_nw              (ready_o_gather_nw[3][6]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[3][6]),
    .data_i_merge_nw                (data_o_merge_nw[3][6]),
    .ready_o_merge_nw               (ready_i_merge_nw[3][6]),
    .valid_o_merge_nw               (valid_i_merge_nw[3][6]),
    .data_o_merge_nw                (data_i_merge_nw[3][6]),
    .ready_i_merge_nw               (ready_o_merge_nw[3][6]),

    .valid_i_cast_pe                (cast_valid_i_3_6),
    .data_i_cast_pe                 (cast_data_i_3_6),
    .ready_o_cast_pe                (cast_ready_o_3_6),
    .valid_o_cast_pe                (cast_valid_o_3_6),
    .data_o_cast_pe                 (cast_data_o_3_6),
    .ready_i_cast_pe                (cast_ready_i_3_6),

    .valid_i_merge_pe               (merge_valid_i_3_6),
    .data_i_merge_pe                (merge_data_i_3_6),
    .ready_o_merge_pe               (merge_ready_o_3_6),
    .valid_o_merge_pe               (merge_valid_o_3_6),
    .data_o_merge_pe                (merge_data_o_3_6),
    .ready_i_merge_pe               (merge_ready_i_3_6),

    .valid_i_gather_pe              (gather_valid_i_3_6),
    .data_i_gather_pe               (gather_data_i_3_6),
    .ready_o_gather_pe              (gather_ready_o_3_6),
    .valid_o_gather_pe              (gather_valid_o_3_6),
    .data_o_gather_pe               (gather_data_o_3_6),
    .ready_i_gather_pe              (gather_ready_i_3_6),

    .credit_upd                     (credit_upd[3][6])
);


network_interface #(
    .cast_out                       (cast_out_3_7),
    .gather_out                     (gather_out_3_7),
    .cast_sid                       (cast_sid_3_7),
    .gather_sid                     (gather_sid_3_7)
)ni_3_7(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[3][7]),
    .data_i_cast_nw                 (data_o_cast_nw[3][7]),
    .ready_o_cast_nw                (ready_i_cast_nw[3][7]),
    .valid_o_cast_nw                (valid_i_cast_nw[3][7]),
    .data_o_cast_nw                 (data_i_cast_nw[3][7]),
    .ready_i_cast_nw                (ready_o_cast_nw[3][7]),

    .valid_i_gather_nw              (valid_o_gather_nw[3][7]),
    .data_i_gather_nw               (data_o_gather_nw[3][7]),
    .ready_o_gather_nw              (ready_i_gather_nw[3][7]),
    .valid_o_gather_nw              (valid_i_gather_nw[3][7]),
    .data_o_gather_nw               (data_i_gather_nw[3][7]),
    .ready_i_gather_nw              (ready_o_gather_nw[3][7]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[3][7]),
    .data_i_merge_nw                (data_o_merge_nw[3][7]),
    .ready_o_merge_nw               (ready_i_merge_nw[3][7]),
    .valid_o_merge_nw               (valid_i_merge_nw[3][7]),
    .data_o_merge_nw                (data_i_merge_nw[3][7]),
    .ready_i_merge_nw               (ready_o_merge_nw[3][7]),

    .valid_i_cast_pe                (cast_valid_i_3_7),
    .data_i_cast_pe                 (cast_data_i_3_7),
    .ready_o_cast_pe                (cast_ready_o_3_7),
    .valid_o_cast_pe                (cast_valid_o_3_7),
    .data_o_cast_pe                 (cast_data_o_3_7),
    .ready_i_cast_pe                (cast_ready_i_3_7),

    .valid_i_merge_pe               (merge_valid_i_3_7),
    .data_i_merge_pe                (merge_data_i_3_7),
    .ready_o_merge_pe               (merge_ready_o_3_7),
    .valid_o_merge_pe               (merge_valid_o_3_7),
    .data_o_merge_pe                (merge_data_o_3_7),
    .ready_i_merge_pe               (merge_ready_i_3_7),

    .valid_i_gather_pe              (gather_valid_i_3_7),
    .data_i_gather_pe               (gather_data_i_3_7),
    .ready_o_gather_pe              (gather_ready_o_3_7),
    .valid_o_gather_pe              (gather_valid_o_3_7),
    .data_o_gather_pe               (gather_data_o_3_7),
    .ready_i_gather_pe              (gather_ready_i_3_7),

    .credit_upd                     (credit_upd[3][7])
);


network_interface #(
    .cast_out                       (cast_out_3_8),
    .gather_out                     (gather_out_3_8),
    .cast_sid                       (cast_sid_3_8),
    .gather_sid                     (gather_sid_3_8)
)ni_3_8(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[3][8]),
    .data_i_cast_nw                 (data_o_cast_nw[3][8]),
    .ready_o_cast_nw                (ready_i_cast_nw[3][8]),
    .valid_o_cast_nw                (valid_i_cast_nw[3][8]),
    .data_o_cast_nw                 (data_i_cast_nw[3][8]),
    .ready_i_cast_nw                (ready_o_cast_nw[3][8]),

    .valid_i_gather_nw              (valid_o_gather_nw[3][8]),
    .data_i_gather_nw               (data_o_gather_nw[3][8]),
    .ready_o_gather_nw              (ready_i_gather_nw[3][8]),
    .valid_o_gather_nw              (valid_i_gather_nw[3][8]),
    .data_o_gather_nw               (data_i_gather_nw[3][8]),
    .ready_i_gather_nw              (ready_o_gather_nw[3][8]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[3][8]),
    .data_i_merge_nw                (data_o_merge_nw[3][8]),
    .ready_o_merge_nw               (ready_i_merge_nw[3][8]),
    .valid_o_merge_nw               (valid_i_merge_nw[3][8]),
    .data_o_merge_nw                (data_i_merge_nw[3][8]),
    .ready_i_merge_nw               (ready_o_merge_nw[3][8]),

    .valid_i_cast_pe                (cast_valid_i_3_8),
    .data_i_cast_pe                 (cast_data_i_3_8),
    .ready_o_cast_pe                (cast_ready_o_3_8),
    .valid_o_cast_pe                (cast_valid_o_3_8),
    .data_o_cast_pe                 (cast_data_o_3_8),
    .ready_i_cast_pe                (cast_ready_i_3_8),

    .valid_i_merge_pe               (merge_valid_i_3_8),
    .data_i_merge_pe                (merge_data_i_3_8),
    .ready_o_merge_pe               (merge_ready_o_3_8),
    .valid_o_merge_pe               (merge_valid_o_3_8),
    .data_o_merge_pe                (merge_data_o_3_8),
    .ready_i_merge_pe               (merge_ready_i_3_8),

    .valid_i_gather_pe              (gather_valid_i_3_8),
    .data_i_gather_pe               (gather_data_i_3_8),
    .ready_o_gather_pe              (gather_ready_o_3_8),
    .valid_o_gather_pe              (gather_valid_o_3_8),
    .data_o_gather_pe               (gather_data_o_3_8),
    .ready_i_gather_pe              (gather_ready_i_3_8),

    .credit_upd                     (credit_upd[3][8])
);


network_interface #(
    .cast_out                       (cast_out_3_9),
    .gather_out                     (gather_out_3_9),
    .cast_sid                       (cast_sid_3_9),
    .gather_sid                     (gather_sid_3_9)
)ni_3_9(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[3][9]),
    .data_i_cast_nw                 (data_o_cast_nw[3][9]),
    .ready_o_cast_nw                (ready_i_cast_nw[3][9]),
    .valid_o_cast_nw                (valid_i_cast_nw[3][9]),
    .data_o_cast_nw                 (data_i_cast_nw[3][9]),
    .ready_i_cast_nw                (ready_o_cast_nw[3][9]),

    .valid_i_gather_nw              (valid_o_gather_nw[3][9]),
    .data_i_gather_nw               (data_o_gather_nw[3][9]),
    .ready_o_gather_nw              (ready_i_gather_nw[3][9]),
    .valid_o_gather_nw              (valid_i_gather_nw[3][9]),
    .data_o_gather_nw               (data_i_gather_nw[3][9]),
    .ready_i_gather_nw              (ready_o_gather_nw[3][9]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[3][9]),
    .data_i_merge_nw                (data_o_merge_nw[3][9]),
    .ready_o_merge_nw               (ready_i_merge_nw[3][9]),
    .valid_o_merge_nw               (valid_i_merge_nw[3][9]),
    .data_o_merge_nw                (data_i_merge_nw[3][9]),
    .ready_i_merge_nw               (ready_o_merge_nw[3][9]),

    .valid_i_cast_pe                (cast_valid_i_3_9),
    .data_i_cast_pe                 (cast_data_i_3_9),
    .ready_o_cast_pe                (cast_ready_o_3_9),
    .valid_o_cast_pe                (cast_valid_o_3_9),
    .data_o_cast_pe                 (cast_data_o_3_9),
    .ready_i_cast_pe                (cast_ready_i_3_9),

    .valid_i_merge_pe               (merge_valid_i_3_9),
    .data_i_merge_pe                (merge_data_i_3_9),
    .ready_o_merge_pe               (merge_ready_o_3_9),
    .valid_o_merge_pe               (merge_valid_o_3_9),
    .data_o_merge_pe                (merge_data_o_3_9),
    .ready_i_merge_pe               (merge_ready_i_3_9),

    .valid_i_gather_pe              (gather_valid_i_3_9),
    .data_i_gather_pe               (gather_data_i_3_9),
    .ready_o_gather_pe              (gather_ready_o_3_9),
    .valid_o_gather_pe              (gather_valid_o_3_9),
    .data_o_gather_pe               (gather_data_o_3_9),
    .ready_i_gather_pe              (gather_ready_i_3_9),

    .credit_upd                     (credit_upd[3][9])
);


network_interface #(
    .cast_out                       (cast_out_4_0),
    .gather_out                     (gather_out_4_0),
    .cast_sid                       (cast_sid_4_0),
    .gather_sid                     (gather_sid_4_0)
)ni_4_0(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[4][0]),
    .data_i_cast_nw                 (data_o_cast_nw[4][0]),
    .ready_o_cast_nw                (ready_i_cast_nw[4][0]),
    .valid_o_cast_nw                (valid_i_cast_nw[4][0]),
    .data_o_cast_nw                 (data_i_cast_nw[4][0]),
    .ready_i_cast_nw                (ready_o_cast_nw[4][0]),

    .valid_i_gather_nw              (valid_o_gather_nw[4][0]),
    .data_i_gather_nw               (data_o_gather_nw[4][0]),
    .ready_o_gather_nw              (ready_i_gather_nw[4][0]),
    .valid_o_gather_nw              (valid_i_gather_nw[4][0]),
    .data_o_gather_nw               (data_i_gather_nw[4][0]),
    .ready_i_gather_nw              (ready_o_gather_nw[4][0]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[4][0]),
    .data_i_merge_nw                (data_o_merge_nw[4][0]),
    .ready_o_merge_nw               (ready_i_merge_nw[4][0]),
    .valid_o_merge_nw               (valid_i_merge_nw[4][0]),
    .data_o_merge_nw                (data_i_merge_nw[4][0]),
    .ready_i_merge_nw               (ready_o_merge_nw[4][0]),

    .valid_i_cast_pe                (cast_valid_i_4_0),
    .data_i_cast_pe                 (cast_data_i_4_0),
    .ready_o_cast_pe                (cast_ready_o_4_0),
    .valid_o_cast_pe                (cast_valid_o_4_0),
    .data_o_cast_pe                 (cast_data_o_4_0),
    .ready_i_cast_pe                (cast_ready_i_4_0),

    .valid_i_merge_pe               (merge_valid_i_4_0),
    .data_i_merge_pe                (merge_data_i_4_0),
    .ready_o_merge_pe               (merge_ready_o_4_0),
    .valid_o_merge_pe               (merge_valid_o_4_0),
    .data_o_merge_pe                (merge_data_o_4_0),
    .ready_i_merge_pe               (merge_ready_i_4_0),

    .valid_i_gather_pe              (gather_valid_i_4_0),
    .data_i_gather_pe               (gather_data_i_4_0),
    .ready_o_gather_pe              (gather_ready_o_4_0),
    .valid_o_gather_pe              (gather_valid_o_4_0),
    .data_o_gather_pe               (gather_data_o_4_0),
    .ready_i_gather_pe              (gather_ready_i_4_0),

    .credit_upd                     (credit_upd[4][0])
);


network_interface #(
    .cast_out                       (cast_out_4_1),
    .gather_out                     (gather_out_4_1),
    .cast_sid                       (cast_sid_4_1),
    .gather_sid                     (gather_sid_4_1)
)ni_4_1(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[4][1]),
    .data_i_cast_nw                 (data_o_cast_nw[4][1]),
    .ready_o_cast_nw                (ready_i_cast_nw[4][1]),
    .valid_o_cast_nw                (valid_i_cast_nw[4][1]),
    .data_o_cast_nw                 (data_i_cast_nw[4][1]),
    .ready_i_cast_nw                (ready_o_cast_nw[4][1]),

    .valid_i_gather_nw              (valid_o_gather_nw[4][1]),
    .data_i_gather_nw               (data_o_gather_nw[4][1]),
    .ready_o_gather_nw              (ready_i_gather_nw[4][1]),
    .valid_o_gather_nw              (valid_i_gather_nw[4][1]),
    .data_o_gather_nw               (data_i_gather_nw[4][1]),
    .ready_i_gather_nw              (ready_o_gather_nw[4][1]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[4][1]),
    .data_i_merge_nw                (data_o_merge_nw[4][1]),
    .ready_o_merge_nw               (ready_i_merge_nw[4][1]),
    .valid_o_merge_nw               (valid_i_merge_nw[4][1]),
    .data_o_merge_nw                (data_i_merge_nw[4][1]),
    .ready_i_merge_nw               (ready_o_merge_nw[4][1]),

    .valid_i_cast_pe                (cast_valid_i_4_1),
    .data_i_cast_pe                 (cast_data_i_4_1),
    .ready_o_cast_pe                (cast_ready_o_4_1),
    .valid_o_cast_pe                (cast_valid_o_4_1),
    .data_o_cast_pe                 (cast_data_o_4_1),
    .ready_i_cast_pe                (cast_ready_i_4_1),

    .valid_i_merge_pe               (merge_valid_i_4_1),
    .data_i_merge_pe                (merge_data_i_4_1),
    .ready_o_merge_pe               (merge_ready_o_4_1),
    .valid_o_merge_pe               (merge_valid_o_4_1),
    .data_o_merge_pe                (merge_data_o_4_1),
    .ready_i_merge_pe               (merge_ready_i_4_1),

    .valid_i_gather_pe              (gather_valid_i_4_1),
    .data_i_gather_pe               (gather_data_i_4_1),
    .ready_o_gather_pe              (gather_ready_o_4_1),
    .valid_o_gather_pe              (gather_valid_o_4_1),
    .data_o_gather_pe               (gather_data_o_4_1),
    .ready_i_gather_pe              (gather_ready_i_4_1),

    .credit_upd                     (credit_upd[4][1])
);


network_interface #(
    .cast_out                       (cast_out_4_2),
    .gather_out                     (gather_out_4_2),
    .cast_sid                       (cast_sid_4_2),
    .gather_sid                     (gather_sid_4_2)
)ni_4_2(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[4][2]),
    .data_i_cast_nw                 (data_o_cast_nw[4][2]),
    .ready_o_cast_nw                (ready_i_cast_nw[4][2]),
    .valid_o_cast_nw                (valid_i_cast_nw[4][2]),
    .data_o_cast_nw                 (data_i_cast_nw[4][2]),
    .ready_i_cast_nw                (ready_o_cast_nw[4][2]),

    .valid_i_gather_nw              (valid_o_gather_nw[4][2]),
    .data_i_gather_nw               (data_o_gather_nw[4][2]),
    .ready_o_gather_nw              (ready_i_gather_nw[4][2]),
    .valid_o_gather_nw              (valid_i_gather_nw[4][2]),
    .data_o_gather_nw               (data_i_gather_nw[4][2]),
    .ready_i_gather_nw              (ready_o_gather_nw[4][2]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[4][2]),
    .data_i_merge_nw                (data_o_merge_nw[4][2]),
    .ready_o_merge_nw               (ready_i_merge_nw[4][2]),
    .valid_o_merge_nw               (valid_i_merge_nw[4][2]),
    .data_o_merge_nw                (data_i_merge_nw[4][2]),
    .ready_i_merge_nw               (ready_o_merge_nw[4][2]),

    .valid_i_cast_pe                (cast_valid_i_4_2),
    .data_i_cast_pe                 (cast_data_i_4_2),
    .ready_o_cast_pe                (cast_ready_o_4_2),
    .valid_o_cast_pe                (cast_valid_o_4_2),
    .data_o_cast_pe                 (cast_data_o_4_2),
    .ready_i_cast_pe                (cast_ready_i_4_2),

    .valid_i_merge_pe               (merge_valid_i_4_2),
    .data_i_merge_pe                (merge_data_i_4_2),
    .ready_o_merge_pe               (merge_ready_o_4_2),
    .valid_o_merge_pe               (merge_valid_o_4_2),
    .data_o_merge_pe                (merge_data_o_4_2),
    .ready_i_merge_pe               (merge_ready_i_4_2),

    .valid_i_gather_pe              (gather_valid_i_4_2),
    .data_i_gather_pe               (gather_data_i_4_2),
    .ready_o_gather_pe              (gather_ready_o_4_2),
    .valid_o_gather_pe              (gather_valid_o_4_2),
    .data_o_gather_pe               (gather_data_o_4_2),
    .ready_i_gather_pe              (gather_ready_i_4_2),

    .credit_upd                     (credit_upd[4][2])
);


network_interface #(
    .cast_out                       (cast_out_4_3),
    .gather_out                     (gather_out_4_3),
    .cast_sid                       (cast_sid_4_3),
    .gather_sid                     (gather_sid_4_3)
)ni_4_3(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[4][3]),
    .data_i_cast_nw                 (data_o_cast_nw[4][3]),
    .ready_o_cast_nw                (ready_i_cast_nw[4][3]),
    .valid_o_cast_nw                (valid_i_cast_nw[4][3]),
    .data_o_cast_nw                 (data_i_cast_nw[4][3]),
    .ready_i_cast_nw                (ready_o_cast_nw[4][3]),

    .valid_i_gather_nw              (valid_o_gather_nw[4][3]),
    .data_i_gather_nw               (data_o_gather_nw[4][3]),
    .ready_o_gather_nw              (ready_i_gather_nw[4][3]),
    .valid_o_gather_nw              (valid_i_gather_nw[4][3]),
    .data_o_gather_nw               (data_i_gather_nw[4][3]),
    .ready_i_gather_nw              (ready_o_gather_nw[4][3]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[4][3]),
    .data_i_merge_nw                (data_o_merge_nw[4][3]),
    .ready_o_merge_nw               (ready_i_merge_nw[4][3]),
    .valid_o_merge_nw               (valid_i_merge_nw[4][3]),
    .data_o_merge_nw                (data_i_merge_nw[4][3]),
    .ready_i_merge_nw               (ready_o_merge_nw[4][3]),

    .valid_i_cast_pe                (cast_valid_i_4_3),
    .data_i_cast_pe                 (cast_data_i_4_3),
    .ready_o_cast_pe                (cast_ready_o_4_3),
    .valid_o_cast_pe                (cast_valid_o_4_3),
    .data_o_cast_pe                 (cast_data_o_4_3),
    .ready_i_cast_pe                (cast_ready_i_4_3),

    .valid_i_merge_pe               (merge_valid_i_4_3),
    .data_i_merge_pe                (merge_data_i_4_3),
    .ready_o_merge_pe               (merge_ready_o_4_3),
    .valid_o_merge_pe               (merge_valid_o_4_3),
    .data_o_merge_pe                (merge_data_o_4_3),
    .ready_i_merge_pe               (merge_ready_i_4_3),

    .valid_i_gather_pe              (gather_valid_i_4_3),
    .data_i_gather_pe               (gather_data_i_4_3),
    .ready_o_gather_pe              (gather_ready_o_4_3),
    .valid_o_gather_pe              (gather_valid_o_4_3),
    .data_o_gather_pe               (gather_data_o_4_3),
    .ready_i_gather_pe              (gather_ready_i_4_3),

    .credit_upd                     (credit_upd[4][3])
);


network_interface #(
    .cast_out                       (cast_out_4_4),
    .gather_out                     (gather_out_4_4),
    .cast_sid                       (cast_sid_4_4),
    .gather_sid                     (gather_sid_4_4)
)ni_4_4(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[4][4]),
    .data_i_cast_nw                 (data_o_cast_nw[4][4]),
    .ready_o_cast_nw                (ready_i_cast_nw[4][4]),
    .valid_o_cast_nw                (valid_i_cast_nw[4][4]),
    .data_o_cast_nw                 (data_i_cast_nw[4][4]),
    .ready_i_cast_nw                (ready_o_cast_nw[4][4]),

    .valid_i_gather_nw              (valid_o_gather_nw[4][4]),
    .data_i_gather_nw               (data_o_gather_nw[4][4]),
    .ready_o_gather_nw              (ready_i_gather_nw[4][4]),
    .valid_o_gather_nw              (valid_i_gather_nw[4][4]),
    .data_o_gather_nw               (data_i_gather_nw[4][4]),
    .ready_i_gather_nw              (ready_o_gather_nw[4][4]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[4][4]),
    .data_i_merge_nw                (data_o_merge_nw[4][4]),
    .ready_o_merge_nw               (ready_i_merge_nw[4][4]),
    .valid_o_merge_nw               (valid_i_merge_nw[4][4]),
    .data_o_merge_nw                (data_i_merge_nw[4][4]),
    .ready_i_merge_nw               (ready_o_merge_nw[4][4]),

    .valid_i_cast_pe                (cast_valid_i_4_4),
    .data_i_cast_pe                 (cast_data_i_4_4),
    .ready_o_cast_pe                (cast_ready_o_4_4),
    .valid_o_cast_pe                (cast_valid_o_4_4),
    .data_o_cast_pe                 (cast_data_o_4_4),
    .ready_i_cast_pe                (cast_ready_i_4_4),

    .valid_i_merge_pe               (merge_valid_i_4_4),
    .data_i_merge_pe                (merge_data_i_4_4),
    .ready_o_merge_pe               (merge_ready_o_4_4),
    .valid_o_merge_pe               (merge_valid_o_4_4),
    .data_o_merge_pe                (merge_data_o_4_4),
    .ready_i_merge_pe               (merge_ready_i_4_4),

    .valid_i_gather_pe              (gather_valid_i_4_4),
    .data_i_gather_pe               (gather_data_i_4_4),
    .ready_o_gather_pe              (gather_ready_o_4_4),
    .valid_o_gather_pe              (gather_valid_o_4_4),
    .data_o_gather_pe               (gather_data_o_4_4),
    .ready_i_gather_pe              (gather_ready_i_4_4),

    .credit_upd                     (credit_upd[4][4])
);


network_interface #(
    .cast_out                       (cast_out_4_5),
    .gather_out                     (gather_out_4_5),
    .cast_sid                       (cast_sid_4_5),
    .gather_sid                     (gather_sid_4_5)
)ni_4_5(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[4][5]),
    .data_i_cast_nw                 (data_o_cast_nw[4][5]),
    .ready_o_cast_nw                (ready_i_cast_nw[4][5]),
    .valid_o_cast_nw                (valid_i_cast_nw[4][5]),
    .data_o_cast_nw                 (data_i_cast_nw[4][5]),
    .ready_i_cast_nw                (ready_o_cast_nw[4][5]),

    .valid_i_gather_nw              (valid_o_gather_nw[4][5]),
    .data_i_gather_nw               (data_o_gather_nw[4][5]),
    .ready_o_gather_nw              (ready_i_gather_nw[4][5]),
    .valid_o_gather_nw              (valid_i_gather_nw[4][5]),
    .data_o_gather_nw               (data_i_gather_nw[4][5]),
    .ready_i_gather_nw              (ready_o_gather_nw[4][5]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[4][5]),
    .data_i_merge_nw                (data_o_merge_nw[4][5]),
    .ready_o_merge_nw               (ready_i_merge_nw[4][5]),
    .valid_o_merge_nw               (valid_i_merge_nw[4][5]),
    .data_o_merge_nw                (data_i_merge_nw[4][5]),
    .ready_i_merge_nw               (ready_o_merge_nw[4][5]),

    .valid_i_cast_pe                (cast_valid_i_4_5),
    .data_i_cast_pe                 (cast_data_i_4_5),
    .ready_o_cast_pe                (cast_ready_o_4_5),
    .valid_o_cast_pe                (cast_valid_o_4_5),
    .data_o_cast_pe                 (cast_data_o_4_5),
    .ready_i_cast_pe                (cast_ready_i_4_5),

    .valid_i_merge_pe               (merge_valid_i_4_5),
    .data_i_merge_pe                (merge_data_i_4_5),
    .ready_o_merge_pe               (merge_ready_o_4_5),
    .valid_o_merge_pe               (merge_valid_o_4_5),
    .data_o_merge_pe                (merge_data_o_4_5),
    .ready_i_merge_pe               (merge_ready_i_4_5),

    .valid_i_gather_pe              (gather_valid_i_4_5),
    .data_i_gather_pe               (gather_data_i_4_5),
    .ready_o_gather_pe              (gather_ready_o_4_5),
    .valid_o_gather_pe              (gather_valid_o_4_5),
    .data_o_gather_pe               (gather_data_o_4_5),
    .ready_i_gather_pe              (gather_ready_i_4_5),

    .credit_upd                     (credit_upd[4][5])
);


network_interface #(
    .cast_out                       (cast_out_4_6),
    .gather_out                     (gather_out_4_6),
    .cast_sid                       (cast_sid_4_6),
    .gather_sid                     (gather_sid_4_6)
)ni_4_6(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[4][6]),
    .data_i_cast_nw                 (data_o_cast_nw[4][6]),
    .ready_o_cast_nw                (ready_i_cast_nw[4][6]),
    .valid_o_cast_nw                (valid_i_cast_nw[4][6]),
    .data_o_cast_nw                 (data_i_cast_nw[4][6]),
    .ready_i_cast_nw                (ready_o_cast_nw[4][6]),

    .valid_i_gather_nw              (valid_o_gather_nw[4][6]),
    .data_i_gather_nw               (data_o_gather_nw[4][6]),
    .ready_o_gather_nw              (ready_i_gather_nw[4][6]),
    .valid_o_gather_nw              (valid_i_gather_nw[4][6]),
    .data_o_gather_nw               (data_i_gather_nw[4][6]),
    .ready_i_gather_nw              (ready_o_gather_nw[4][6]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[4][6]),
    .data_i_merge_nw                (data_o_merge_nw[4][6]),
    .ready_o_merge_nw               (ready_i_merge_nw[4][6]),
    .valid_o_merge_nw               (valid_i_merge_nw[4][6]),
    .data_o_merge_nw                (data_i_merge_nw[4][6]),
    .ready_i_merge_nw               (ready_o_merge_nw[4][6]),

    .valid_i_cast_pe                (cast_valid_i_4_6),
    .data_i_cast_pe                 (cast_data_i_4_6),
    .ready_o_cast_pe                (cast_ready_o_4_6),
    .valid_o_cast_pe                (cast_valid_o_4_6),
    .data_o_cast_pe                 (cast_data_o_4_6),
    .ready_i_cast_pe                (cast_ready_i_4_6),

    .valid_i_merge_pe               (merge_valid_i_4_6),
    .data_i_merge_pe                (merge_data_i_4_6),
    .ready_o_merge_pe               (merge_ready_o_4_6),
    .valid_o_merge_pe               (merge_valid_o_4_6),
    .data_o_merge_pe                (merge_data_o_4_6),
    .ready_i_merge_pe               (merge_ready_i_4_6),

    .valid_i_gather_pe              (gather_valid_i_4_6),
    .data_i_gather_pe               (gather_data_i_4_6),
    .ready_o_gather_pe              (gather_ready_o_4_6),
    .valid_o_gather_pe              (gather_valid_o_4_6),
    .data_o_gather_pe               (gather_data_o_4_6),
    .ready_i_gather_pe              (gather_ready_i_4_6),

    .credit_upd                     (credit_upd[4][6])
);


network_interface #(
    .cast_out                       (cast_out_4_7),
    .gather_out                     (gather_out_4_7),
    .cast_sid                       (cast_sid_4_7),
    .gather_sid                     (gather_sid_4_7)
)ni_4_7(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[4][7]),
    .data_i_cast_nw                 (data_o_cast_nw[4][7]),
    .ready_o_cast_nw                (ready_i_cast_nw[4][7]),
    .valid_o_cast_nw                (valid_i_cast_nw[4][7]),
    .data_o_cast_nw                 (data_i_cast_nw[4][7]),
    .ready_i_cast_nw                (ready_o_cast_nw[4][7]),

    .valid_i_gather_nw              (valid_o_gather_nw[4][7]),
    .data_i_gather_nw               (data_o_gather_nw[4][7]),
    .ready_o_gather_nw              (ready_i_gather_nw[4][7]),
    .valid_o_gather_nw              (valid_i_gather_nw[4][7]),
    .data_o_gather_nw               (data_i_gather_nw[4][7]),
    .ready_i_gather_nw              (ready_o_gather_nw[4][7]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[4][7]),
    .data_i_merge_nw                (data_o_merge_nw[4][7]),
    .ready_o_merge_nw               (ready_i_merge_nw[4][7]),
    .valid_o_merge_nw               (valid_i_merge_nw[4][7]),
    .data_o_merge_nw                (data_i_merge_nw[4][7]),
    .ready_i_merge_nw               (ready_o_merge_nw[4][7]),

    .valid_i_cast_pe                (cast_valid_i_4_7),
    .data_i_cast_pe                 (cast_data_i_4_7),
    .ready_o_cast_pe                (cast_ready_o_4_7),
    .valid_o_cast_pe                (cast_valid_o_4_7),
    .data_o_cast_pe                 (cast_data_o_4_7),
    .ready_i_cast_pe                (cast_ready_i_4_7),

    .valid_i_merge_pe               (merge_valid_i_4_7),
    .data_i_merge_pe                (merge_data_i_4_7),
    .ready_o_merge_pe               (merge_ready_o_4_7),
    .valid_o_merge_pe               (merge_valid_o_4_7),
    .data_o_merge_pe                (merge_data_o_4_7),
    .ready_i_merge_pe               (merge_ready_i_4_7),

    .valid_i_gather_pe              (gather_valid_i_4_7),
    .data_i_gather_pe               (gather_data_i_4_7),
    .ready_o_gather_pe              (gather_ready_o_4_7),
    .valid_o_gather_pe              (gather_valid_o_4_7),
    .data_o_gather_pe               (gather_data_o_4_7),
    .ready_i_gather_pe              (gather_ready_i_4_7),

    .credit_upd                     (credit_upd[4][7])
);


network_interface #(
    .cast_out                       (cast_out_4_8),
    .gather_out                     (gather_out_4_8),
    .cast_sid                       (cast_sid_4_8),
    .gather_sid                     (gather_sid_4_8)
)ni_4_8(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[4][8]),
    .data_i_cast_nw                 (data_o_cast_nw[4][8]),
    .ready_o_cast_nw                (ready_i_cast_nw[4][8]),
    .valid_o_cast_nw                (valid_i_cast_nw[4][8]),
    .data_o_cast_nw                 (data_i_cast_nw[4][8]),
    .ready_i_cast_nw                (ready_o_cast_nw[4][8]),

    .valid_i_gather_nw              (valid_o_gather_nw[4][8]),
    .data_i_gather_nw               (data_o_gather_nw[4][8]),
    .ready_o_gather_nw              (ready_i_gather_nw[4][8]),
    .valid_o_gather_nw              (valid_i_gather_nw[4][8]),
    .data_o_gather_nw               (data_i_gather_nw[4][8]),
    .ready_i_gather_nw              (ready_o_gather_nw[4][8]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[4][8]),
    .data_i_merge_nw                (data_o_merge_nw[4][8]),
    .ready_o_merge_nw               (ready_i_merge_nw[4][8]),
    .valid_o_merge_nw               (valid_i_merge_nw[4][8]),
    .data_o_merge_nw                (data_i_merge_nw[4][8]),
    .ready_i_merge_nw               (ready_o_merge_nw[4][8]),

    .valid_i_cast_pe                (cast_valid_i_4_8),
    .data_i_cast_pe                 (cast_data_i_4_8),
    .ready_o_cast_pe                (cast_ready_o_4_8),
    .valid_o_cast_pe                (cast_valid_o_4_8),
    .data_o_cast_pe                 (cast_data_o_4_8),
    .ready_i_cast_pe                (cast_ready_i_4_8),

    .valid_i_merge_pe               (merge_valid_i_4_8),
    .data_i_merge_pe                (merge_data_i_4_8),
    .ready_o_merge_pe               (merge_ready_o_4_8),
    .valid_o_merge_pe               (merge_valid_o_4_8),
    .data_o_merge_pe                (merge_data_o_4_8),
    .ready_i_merge_pe               (merge_ready_i_4_8),

    .valid_i_gather_pe              (gather_valid_i_4_8),
    .data_i_gather_pe               (gather_data_i_4_8),
    .ready_o_gather_pe              (gather_ready_o_4_8),
    .valid_o_gather_pe              (gather_valid_o_4_8),
    .data_o_gather_pe               (gather_data_o_4_8),
    .ready_i_gather_pe              (gather_ready_i_4_8),

    .credit_upd                     (credit_upd[4][8])
);


network_interface #(
    .cast_out                       (cast_out_4_9),
    .gather_out                     (gather_out_4_9),
    .cast_sid                       (cast_sid_4_9),
    .gather_sid                     (gather_sid_4_9)
)ni_4_9(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[4][9]),
    .data_i_cast_nw                 (data_o_cast_nw[4][9]),
    .ready_o_cast_nw                (ready_i_cast_nw[4][9]),
    .valid_o_cast_nw                (valid_i_cast_nw[4][9]),
    .data_o_cast_nw                 (data_i_cast_nw[4][9]),
    .ready_i_cast_nw                (ready_o_cast_nw[4][9]),

    .valid_i_gather_nw              (valid_o_gather_nw[4][9]),
    .data_i_gather_nw               (data_o_gather_nw[4][9]),
    .ready_o_gather_nw              (ready_i_gather_nw[4][9]),
    .valid_o_gather_nw              (valid_i_gather_nw[4][9]),
    .data_o_gather_nw               (data_i_gather_nw[4][9]),
    .ready_i_gather_nw              (ready_o_gather_nw[4][9]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[4][9]),
    .data_i_merge_nw                (data_o_merge_nw[4][9]),
    .ready_o_merge_nw               (ready_i_merge_nw[4][9]),
    .valid_o_merge_nw               (valid_i_merge_nw[4][9]),
    .data_o_merge_nw                (data_i_merge_nw[4][9]),
    .ready_i_merge_nw               (ready_o_merge_nw[4][9]),

    .valid_i_cast_pe                (cast_valid_i_4_9),
    .data_i_cast_pe                 (cast_data_i_4_9),
    .ready_o_cast_pe                (cast_ready_o_4_9),
    .valid_o_cast_pe                (cast_valid_o_4_9),
    .data_o_cast_pe                 (cast_data_o_4_9),
    .ready_i_cast_pe                (cast_ready_i_4_9),

    .valid_i_merge_pe               (merge_valid_i_4_9),
    .data_i_merge_pe                (merge_data_i_4_9),
    .ready_o_merge_pe               (merge_ready_o_4_9),
    .valid_o_merge_pe               (merge_valid_o_4_9),
    .data_o_merge_pe                (merge_data_o_4_9),
    .ready_i_merge_pe               (merge_ready_i_4_9),

    .valid_i_gather_pe              (gather_valid_i_4_9),
    .data_i_gather_pe               (gather_data_i_4_9),
    .ready_o_gather_pe              (gather_ready_o_4_9),
    .valid_o_gather_pe              (gather_valid_o_4_9),
    .data_o_gather_pe               (gather_data_o_4_9),
    .ready_i_gather_pe              (gather_ready_i_4_9),

    .credit_upd                     (credit_upd[4][9])
);

endmodule
