localparam isUBM_list_0_0[`CN] = '{0,0,0,0,0};
localparam isUBM_list_0_1[`CN] = '{0,0,0,0,0};
localparam isUBM_list_0_2[`CN] = '{0,0,0,0,0};
localparam isUBM_list_0_3[`CN] = '{0,0,0,0,0};
localparam isUBM_list_0_4[`CN] = '{0,0,0,0,0};
localparam isUBM_list_0_5[`CN] = '{0,0,0,0,0};
localparam isUBM_list_0_6[`CN] = '{0,0,0,0,0};
localparam isUBM_list_0_7[`CN] = '{0,0,0,0,0};
localparam isUBM_list_0_8[`CN] = '{0,0,0,0,0};
localparam isUBM_list_0_9[`CN] = '{0,0,0,0,0};
localparam isUBM_list_0_10[`CN] = '{0,0,0,0,0};
localparam isUBM_list_1_0[`CN] = '{0,0,0,0,0};
localparam isUBM_list_1_1[`CN] = '{0,0,0,0,0};
localparam isUBM_list_1_2[`CN] = '{0,0,0,0,0};
localparam isUBM_list_1_3[`CN] = '{0,0,0,0,0};
localparam isUBM_list_1_4[`CN] = '{0,0,0,0,0};
localparam isUBM_list_1_5[`CN] = '{0,0,0,0,0};
localparam isUBM_list_1_6[`CN] = '{0,0,0,0,0};
localparam isUBM_list_1_7[`CN] = '{0,0,0,0,0};
localparam isUBM_list_1_8[`CN] = '{0,0,0,0,0};
localparam isUBM_list_1_9[`CN] = '{0,0,0,0,0};
localparam isUBM_list_1_10[`CN] = '{0,0,0,0,0};
localparam isUBM_list_2_0[`CN] = '{0,0,0,0,0};
localparam isUBM_list_2_1[`CN] = '{0,0,0,0,0};
localparam isUBM_list_2_2[`CN] = '{0,0,0,0,0};
localparam isUBM_list_2_3[`CN] = '{0,0,0,0,0};
localparam isUBM_list_2_4[`CN] = '{0,0,0,0,0};
localparam isUBM_list_2_5[`CN] = '{0,0,0,0,0};
localparam isUBM_list_2_6[`CN] = '{0,0,0,0,0};
localparam isUBM_list_2_7[`CN] = '{0,0,0,0,0};
localparam isUBM_list_2_8[`CN] = '{0,0,0,0,0};
localparam isUBM_list_2_9[`CN] = '{0,0,0,0,0};
localparam isUBM_list_2_10[`CN] = '{0,0,0,0,0};
localparam isUBM_list_3_0[`CN] = '{0,0,0,0,0};
localparam isUBM_list_3_1[`CN] = '{0,0,0,0,0};
localparam isUBM_list_3_2[`CN] = '{0,0,0,0,0};
localparam isUBM_list_3_3[`CN] = '{0,0,0,0,0};
localparam isUBM_list_3_4[`CN] = '{0,0,0,0,0};
localparam isUBM_list_3_5[`CN] = '{0,0,0,0,0};
localparam isUBM_list_3_6[`CN] = '{0,0,0,0,0};
localparam isUBM_list_3_7[`CN] = '{0,0,0,0,0};
localparam isUBM_list_3_8[`CN] = '{0,0,0,0,0};
localparam isUBM_list_3_9[`CN] = '{0,0,0,0,0};
localparam isUBM_list_3_10[`CN] = '{0,0,0,0,0};
localparam isUBM_list_4_0[`CN] = '{0,0,0,0,0};
localparam isUBM_list_4_1[`CN] = '{0,0,0,0,0};
localparam isUBM_list_4_2[`CN] = '{0,0,0,0,0};
localparam isUBM_list_4_3[`CN] = '{0,0,0,0,0};
localparam isUBM_list_4_4[`CN] = '{0,0,0,0,0};
localparam isUBM_list_4_5[`CN] = '{0,0,0,0,0};
localparam isUBM_list_4_6[`CN] = '{0,0,0,0,0};
localparam isUBM_list_4_7[`CN] = '{0,0,0,0,0};
localparam isUBM_list_4_8[`CN] = '{0,0,0,0,0};
localparam isUBM_list_4_9[`CN] = '{0,0,0,0,0};
localparam isUBM_list_4_10[`CN] = '{0,0,0,0,0};
localparam isFC_list_0_0[`CN] = '{0,0,0,0,0};
localparam isFC_list_0_1[`CN] = '{0,0,0,0,0};
localparam isFC_list_0_2[`CN] = '{1,0,0,0,0};
localparam isFC_list_0_3[`CN] = '{0,0,0,0,0};
localparam isFC_list_0_4[`CN] = '{1,0,0,0,0};
localparam isFC_list_0_5[`CN] = '{0,0,0,0,0};
localparam isFC_list_0_6[`CN] = '{1,0,0,0,0};
localparam isFC_list_0_7[`CN] = '{0,0,0,0,0};
localparam isFC_list_0_8[`CN] = '{1,0,0,0,0};
localparam isFC_list_0_9[`CN] = '{0,0,0,0,0};
localparam isFC_list_0_10[`CN] = '{0,0,0,0,0};
localparam isFC_list_1_0[`CN] = '{0,0,0,0,0};
localparam isFC_list_1_1[`CN] = '{0,0,0,0,0};
localparam isFC_list_1_2[`CN] = '{0,0,0,0,0};
localparam isFC_list_1_3[`CN] = '{0,0,0,0,0};
localparam isFC_list_1_4[`CN] = '{1,0,0,0,0};
localparam isFC_list_1_5[`CN] = '{0,0,0,0,0};
localparam isFC_list_1_6[`CN] = '{0,0,0,0,0};
localparam isFC_list_1_7[`CN] = '{0,0,0,0,0};
localparam isFC_list_1_8[`CN] = '{0,0,0,0,0};
localparam isFC_list_1_9[`CN] = '{0,0,0,0,0};
localparam isFC_list_1_10[`CN] = '{0,0,0,0,0};
localparam isFC_list_2_0[`CN] = '{0,0,0,0,0};
localparam isFC_list_2_1[`CN] = '{0,0,0,0,0};
localparam isFC_list_2_2[`CN] = '{1,0,0,0,0};
localparam isFC_list_2_3[`CN] = '{0,0,0,0,0};
localparam isFC_list_2_4[`CN] = '{0,0,0,0,0};
localparam isFC_list_2_5[`CN] = '{1,0,0,0,0};
localparam isFC_list_2_6[`CN] = '{0,0,0,0,0};
localparam isFC_list_2_7[`CN] = '{0,0,0,0,0};
localparam isFC_list_2_8[`CN] = '{0,0,0,0,0};
localparam isFC_list_2_9[`CN] = '{0,0,0,0,0};
localparam isFC_list_2_10[`CN] = '{0,0,0,0,0};
localparam isFC_list_3_0[`CN] = '{0,0,0,0,0};
localparam isFC_list_3_1[`CN] = '{0,0,0,0,0};
localparam isFC_list_3_2[`CN] = '{0,0,0,0,0};
localparam isFC_list_3_3[`CN] = '{0,0,0,0,0};
localparam isFC_list_3_4[`CN] = '{0,0,0,0,0};
localparam isFC_list_3_5[`CN] = '{0,0,0,0,0};
localparam isFC_list_3_6[`CN] = '{0,0,0,0,0};
localparam isFC_list_3_7[`CN] = '{0,0,0,0,0};
localparam isFC_list_3_8[`CN] = '{1,0,0,0,0};
localparam isFC_list_3_9[`CN] = '{0,0,0,0,0};
localparam isFC_list_3_10[`CN] = '{0,0,0,0,0};
localparam isFC_list_4_0[`CN] = '{0,0,0,0,0};
localparam isFC_list_4_1[`CN] = '{0,0,0,0,0};
localparam isFC_list_4_2[`CN] = '{0,0,0,0,0};
localparam isFC_list_4_3[`CN] = '{0,0,0,0,0};
localparam isFC_list_4_4[`CN] = '{0,0,0,0,0};
localparam isFC_list_4_5[`CN] = '{0,0,0,0,0};
localparam isFC_list_4_6[`CN] = '{0,0,0,0,0};
localparam isFC_list_4_7[`CN] = '{0,0,0,0,0};
localparam isFC_list_4_8[`CN] = '{0,0,0,0,0};
localparam isFC_list_4_9[`CN] = '{0,0,0,0,0};
localparam isFC_list_4_10[`CN] = '{0,0,0,0,0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_0_0[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_0_1[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_0_2[`CN] = '{55'b0000000000000000000000000000000000111100000000000000000,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_0_3[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_0_4[`CN] = '{55'b0000000000000000000000000001101010000000000000000000000,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_0_5[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_0_6[`CN] = '{55'b0000000000100110010000000000000000000000000000000000000,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_0_7[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_0_8[`CN] = '{55'b0001001101000000000000000000000000000000000000000000000,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_0_9[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_0_10[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_1_0[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_1_1[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_1_2[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_1_3[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_1_4[`CN] = '{55'b0000000000000000100010010000010000000000000000000000000,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_1_5[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_1_6[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_1_7[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_1_8[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_1_9[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_1_10[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_2_0[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_2_1[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_2_2[`CN] = '{55'b0000000000000000000000000000000000000011110000000000000,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_2_3[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_2_4[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_2_5[`CN] = '{55'b0000000000000001000001101000000000000000000000000000000,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_2_6[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_2_7[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_2_8[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_2_9[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_2_10[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_3_0[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_3_1[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_3_2[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_3_3[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_3_4[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_3_5[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_3_6[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_3_7[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_3_8[`CN] = '{55'b0010110010000000000000000000000000000000000000000000000,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_3_9[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_3_10[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_4_0[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_4_1[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_4_2[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_4_3[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_4_4[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_4_5[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_4_6[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_4_7[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_4_8[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_4_9[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_4_10[`CN] = '{55'b0,55'b0,55'b0,55'b0,55'b0};
localparam int FCpl_list_0_0[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_0_1[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_0_2[`CN] = '{`PKT_LEN,0,0,0,0};
localparam int FCpl_list_0_3[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_0_4[`CN] = '{`PKT_LEN,0,0,0,0};
localparam int FCpl_list_0_5[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_0_6[`CN] = '{`PKT_LEN,0,0,0,0};
localparam int FCpl_list_0_7[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_0_8[`CN] = '{`PKT_LEN,0,0,0,0};
localparam int FCpl_list_0_9[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_0_10[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_1_0[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_1_1[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_1_2[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_1_3[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_1_4[`CN] = '{`PKT_LEN,0,0,0,0};
localparam int FCpl_list_1_5[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_1_6[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_1_7[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_1_8[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_1_9[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_1_10[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_2_0[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_2_1[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_2_2[`CN] = '{`PKT_LEN,0,0,0,0};
localparam int FCpl_list_2_3[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_2_4[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_2_5[`CN] = '{`PKT_LEN,0,0,0,0};
localparam int FCpl_list_2_6[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_2_7[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_2_8[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_2_9[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_2_10[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_3_0[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_3_1[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_3_2[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_3_3[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_3_4[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_3_5[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_3_6[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_3_7[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_3_8[`CN] = '{`PKT_LEN,0,0,0,0};
localparam int FCpl_list_3_9[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_3_10[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_4_0[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_4_1[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_4_2[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_4_3[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_4_4[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_4_5[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_4_6[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_4_7[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_4_8[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_4_9[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_4_10[`CN] = '{0,0,0,0,0};
localparam string rt_file_list_0_0[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_0_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_0_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_0_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_0_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_0_4"};
localparam string rt_file_list_0_1[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_1_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_1_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_1_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_1_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_1_4"};
localparam string rt_file_list_0_2[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_2_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_2_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_2_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_2_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_2_4"};
localparam string rt_file_list_0_3[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_3_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_3_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_3_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_3_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_3_4"};
localparam string rt_file_list_0_4[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_4_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_4_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_4_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_4_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_4_4"};
localparam string rt_file_list_0_5[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_5_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_5_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_5_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_5_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_5_4"};
localparam string rt_file_list_0_6[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_6_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_6_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_6_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_6_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_6_4"};
localparam string rt_file_list_0_7[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_7_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_7_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_7_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_7_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_7_4"};
localparam string rt_file_list_0_8[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_8_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_8_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_8_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_8_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_8_4"};
localparam string rt_file_list_0_9[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_9_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_9_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_9_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_9_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_9_4"};
localparam string rt_file_list_0_10[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_10_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_10_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_10_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_10_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_0_10_4"};
localparam string rt_file_list_1_0[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_0_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_0_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_0_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_0_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_0_4"};
localparam string rt_file_list_1_1[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_1_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_1_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_1_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_1_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_1_4"};
localparam string rt_file_list_1_2[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_2_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_2_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_2_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_2_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_2_4"};
localparam string rt_file_list_1_3[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_3_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_3_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_3_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_3_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_3_4"};
localparam string rt_file_list_1_4[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_4_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_4_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_4_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_4_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_4_4"};
localparam string rt_file_list_1_5[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_5_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_5_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_5_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_5_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_5_4"};
localparam string rt_file_list_1_6[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_6_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_6_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_6_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_6_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_6_4"};
localparam string rt_file_list_1_7[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_7_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_7_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_7_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_7_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_7_4"};
localparam string rt_file_list_1_8[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_8_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_8_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_8_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_8_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_8_4"};
localparam string rt_file_list_1_9[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_9_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_9_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_9_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_9_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_9_4"};
localparam string rt_file_list_1_10[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_10_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_10_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_10_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_10_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_1_10_4"};
localparam string rt_file_list_2_0[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_0_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_0_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_0_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_0_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_0_4"};
localparam string rt_file_list_2_1[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_1_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_1_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_1_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_1_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_1_4"};
localparam string rt_file_list_2_2[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_2_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_2_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_2_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_2_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_2_4"};
localparam string rt_file_list_2_3[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_3_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_3_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_3_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_3_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_3_4"};
localparam string rt_file_list_2_4[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_4_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_4_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_4_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_4_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_4_4"};
localparam string rt_file_list_2_5[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_5_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_5_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_5_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_5_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_5_4"};
localparam string rt_file_list_2_6[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_6_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_6_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_6_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_6_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_6_4"};
localparam string rt_file_list_2_7[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_7_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_7_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_7_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_7_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_7_4"};
localparam string rt_file_list_2_8[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_8_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_8_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_8_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_8_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_8_4"};
localparam string rt_file_list_2_9[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_9_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_9_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_9_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_9_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_9_4"};
localparam string rt_file_list_2_10[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_10_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_10_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_10_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_10_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_2_10_4"};
localparam string rt_file_list_3_0[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_0_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_0_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_0_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_0_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_0_4"};
localparam string rt_file_list_3_1[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_1_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_1_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_1_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_1_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_1_4"};
localparam string rt_file_list_3_2[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_2_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_2_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_2_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_2_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_2_4"};
localparam string rt_file_list_3_3[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_3_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_3_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_3_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_3_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_3_4"};
localparam string rt_file_list_3_4[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_4_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_4_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_4_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_4_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_4_4"};
localparam string rt_file_list_3_5[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_5_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_5_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_5_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_5_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_5_4"};
localparam string rt_file_list_3_6[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_6_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_6_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_6_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_6_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_6_4"};
localparam string rt_file_list_3_7[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_7_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_7_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_7_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_7_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_7_4"};
localparam string rt_file_list_3_8[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_8_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_8_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_8_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_8_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_8_4"};
localparam string rt_file_list_3_9[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_9_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_9_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_9_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_9_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_9_4"};
localparam string rt_file_list_3_10[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_10_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_10_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_10_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_10_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_3_10_4"};
localparam string rt_file_list_4_0[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_0_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_0_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_0_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_0_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_0_4"};
localparam string rt_file_list_4_1[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_1_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_1_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_1_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_1_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_1_4"};
localparam string rt_file_list_4_2[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_2_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_2_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_2_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_2_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_2_4"};
localparam string rt_file_list_4_3[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_3_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_3_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_3_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_3_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_3_4"};
localparam string rt_file_list_4_4[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_4_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_4_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_4_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_4_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_4_4"};
localparam string rt_file_list_4_5[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_5_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_5_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_5_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_5_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_5_4"};
localparam string rt_file_list_4_6[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_6_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_6_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_6_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_6_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_6_4"};
localparam string rt_file_list_4_7[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_7_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_7_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_7_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_7_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_7_4"};
localparam string rt_file_list_4_8[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_8_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_8_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_8_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_8_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_8_4"};
localparam string rt_file_list_4_9[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_9_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_9_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_9_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_9_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_9_4"};
localparam string rt_file_list_4_10[`CN] = '{"/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_10_0","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_10_1","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_10_2","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_10_3","/mnt/c/git/nvcim-comm/behavior_model/test_auto/config/cast_rt_4_10_4"};

