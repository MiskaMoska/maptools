`include "params.svh"
`include "network_config.svh"

module system (
    input       wire                            clk,
    input       wire                            rstn,

    input       wire        [`DW-1:0]           data_i_stab,
    input       wire                            valid_i_stab,
    output      wire                            ready_o_stab,

    output      wire        [`DW-1:0]           data_o_flee0,
    output      wire                            valid_o_flee0,
    input       wire                            ready_i_flee0,
    output      wire        [`DW-1:0]           data_o_flee1,
    output      wire                            valid_o_flee1,
    input       wire                            ready_i_flee1
);

wire [`DW-1:0] cast_data_pe_2_nw[`NOC_WIDTH][`NOC_HEIGHT], merge_data_pe_2_nw[`NOC_WIDTH][`NOC_HEIGHT], gather_data_pe_2_nw[`NOC_WIDTH][`NOC_HEIGHT], cast_data_nw_2_pe[`NOC_WIDTH][`NOC_HEIGHT], merge_data_nw_2_pe[`NOC_WIDTH][`NOC_HEIGHT], gather_data_nw_2_pe[`NOC_WIDTH][`NOC_HEIGHT];
wire  cast_valid_pe_2_nw[`NOC_WIDTH][`NOC_HEIGHT], merge_valid_pe_2_nw[`NOC_WIDTH][`NOC_HEIGHT], gather_valid_pe_2_nw[`NOC_WIDTH][`NOC_HEIGHT], cast_valid_nw_2_pe[`NOC_WIDTH][`NOC_HEIGHT], merge_valid_nw_2_pe[`NOC_WIDTH][`NOC_HEIGHT], gather_valid_nw_2_pe[`NOC_WIDTH][`NOC_HEIGHT];
wire  cast_ready_pe_2_nw[`NOC_WIDTH][`NOC_HEIGHT], merge_ready_pe_2_nw[`NOC_WIDTH][`NOC_HEIGHT], gather_ready_pe_2_nw[`NOC_WIDTH][`NOC_HEIGHT], cast_ready_nw_2_pe[`NOC_WIDTH][`NOC_HEIGHT], merge_ready_nw_2_pe[`NOC_WIDTH][`NOC_HEIGHT], gather_ready_nw_2_pe[`NOC_WIDTH][`NOC_HEIGHT];

network nw(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .data_i_stab                                       (data_i_stab),
    .valid_i_stab                                      (valid_i_stab),
    .ready_o_stab                                      (ready_o_stab),
    .data_o_flee0                                      (data_o_flee0),
    .valid_o_flee0                                     (valid_o_flee0),
    .ready_i_flee0                                     (ready_i_flee0),
    .data_o_flee1                                      (data_o_flee1),
    .valid_o_flee1                                     (valid_o_flee1),
    .ready_i_flee1                                     (ready_i_flee1),

    .cast_data_i_0_0                               (cast_data_pe_2_nw[0][0]),
    .cast_valid_i_0_0                              (cast_valid_pe_2_nw[0][0]),
    .cast_ready_o_0_0                              (cast_ready_nw_2_pe[0][0]),
    .merge_data_i_0_0                              (merge_data_pe_2_nw[0][0]),
    .merge_valid_i_0_0                             (merge_valid_pe_2_nw[0][0]),
    .merge_ready_o_0_0                             (merge_ready_nw_2_pe[0][0]),
    .gather_data_i_0_0                             (gather_data_pe_2_nw[0][0]),
    .gather_valid_i_0_0                            (gather_valid_pe_2_nw[0][0]),
    .gather_ready_o_0_0                            (gather_ready_nw_2_pe[0][0]),

    .cast_data_o_0_0                               (cast_data_nw_2_pe[0][0]),
    .cast_valid_o_0_0                              (cast_valid_nw_2_pe[0][0]),
    .cast_ready_i_0_0                              (cast_ready_pe_2_nw[0][0]),
    .merge_data_o_0_0                              (merge_data_nw_2_pe[0][0]),
    .merge_valid_o_0_0                             (merge_valid_nw_2_pe[0][0]),
    .merge_ready_i_0_0                             (merge_ready_pe_2_nw[0][0]),
    .gather_data_o_0_0                             (gather_data_nw_2_pe[0][0]),
    .gather_valid_o_0_0                            (gather_valid_nw_2_pe[0][0]),
    .gather_ready_i_0_0                            (gather_ready_pe_2_nw[0][0]),
    .cast_data_i_0_1                               (cast_data_pe_2_nw[0][1]),
    .cast_valid_i_0_1                              (cast_valid_pe_2_nw[0][1]),
    .cast_ready_o_0_1                              (cast_ready_nw_2_pe[0][1]),
    .merge_data_i_0_1                              (merge_data_pe_2_nw[0][1]),
    .merge_valid_i_0_1                             (merge_valid_pe_2_nw[0][1]),
    .merge_ready_o_0_1                             (merge_ready_nw_2_pe[0][1]),
    .gather_data_i_0_1                             (gather_data_pe_2_nw[0][1]),
    .gather_valid_i_0_1                            (gather_valid_pe_2_nw[0][1]),
    .gather_ready_o_0_1                            (gather_ready_nw_2_pe[0][1]),

    .cast_data_o_0_1                               (cast_data_nw_2_pe[0][1]),
    .cast_valid_o_0_1                              (cast_valid_nw_2_pe[0][1]),
    .cast_ready_i_0_1                              (cast_ready_pe_2_nw[0][1]),
    .merge_data_o_0_1                              (merge_data_nw_2_pe[0][1]),
    .merge_valid_o_0_1                             (merge_valid_nw_2_pe[0][1]),
    .merge_ready_i_0_1                             (merge_ready_pe_2_nw[0][1]),
    .gather_data_o_0_1                             (gather_data_nw_2_pe[0][1]),
    .gather_valid_o_0_1                            (gather_valid_nw_2_pe[0][1]),
    .gather_ready_i_0_1                            (gather_ready_pe_2_nw[0][1]),
    .cast_data_i_0_2                               (cast_data_pe_2_nw[0][2]),
    .cast_valid_i_0_2                              (cast_valid_pe_2_nw[0][2]),
    .cast_ready_o_0_2                              (cast_ready_nw_2_pe[0][2]),
    .merge_data_i_0_2                              (merge_data_pe_2_nw[0][2]),
    .merge_valid_i_0_2                             (merge_valid_pe_2_nw[0][2]),
    .merge_ready_o_0_2                             (merge_ready_nw_2_pe[0][2]),
    .gather_data_i_0_2                             (gather_data_pe_2_nw[0][2]),
    .gather_valid_i_0_2                            (gather_valid_pe_2_nw[0][2]),
    .gather_ready_o_0_2                            (gather_ready_nw_2_pe[0][2]),

    .cast_data_o_0_2                               (cast_data_nw_2_pe[0][2]),
    .cast_valid_o_0_2                              (cast_valid_nw_2_pe[0][2]),
    .cast_ready_i_0_2                              (cast_ready_pe_2_nw[0][2]),
    .merge_data_o_0_2                              (merge_data_nw_2_pe[0][2]),
    .merge_valid_o_0_2                             (merge_valid_nw_2_pe[0][2]),
    .merge_ready_i_0_2                             (merge_ready_pe_2_nw[0][2]),
    .gather_data_o_0_2                             (gather_data_nw_2_pe[0][2]),
    .gather_valid_o_0_2                            (gather_valid_nw_2_pe[0][2]),
    .gather_ready_i_0_2                            (gather_ready_pe_2_nw[0][2]),
    .cast_data_i_0_3                               (cast_data_pe_2_nw[0][3]),
    .cast_valid_i_0_3                              (cast_valid_pe_2_nw[0][3]),
    .cast_ready_o_0_3                              (cast_ready_nw_2_pe[0][3]),
    .merge_data_i_0_3                              (merge_data_pe_2_nw[0][3]),
    .merge_valid_i_0_3                             (merge_valid_pe_2_nw[0][3]),
    .merge_ready_o_0_3                             (merge_ready_nw_2_pe[0][3]),
    .gather_data_i_0_3                             (gather_data_pe_2_nw[0][3]),
    .gather_valid_i_0_3                            (gather_valid_pe_2_nw[0][3]),
    .gather_ready_o_0_3                            (gather_ready_nw_2_pe[0][3]),

    .cast_data_o_0_3                               (cast_data_nw_2_pe[0][3]),
    .cast_valid_o_0_3                              (cast_valid_nw_2_pe[0][3]),
    .cast_ready_i_0_3                              (cast_ready_pe_2_nw[0][3]),
    .merge_data_o_0_3                              (merge_data_nw_2_pe[0][3]),
    .merge_valid_o_0_3                             (merge_valid_nw_2_pe[0][3]),
    .merge_ready_i_0_3                             (merge_ready_pe_2_nw[0][3]),
    .gather_data_o_0_3                             (gather_data_nw_2_pe[0][3]),
    .gather_valid_o_0_3                            (gather_valid_nw_2_pe[0][3]),
    .gather_ready_i_0_3                            (gather_ready_pe_2_nw[0][3]),
    .cast_data_i_0_4                               (cast_data_pe_2_nw[0][4]),
    .cast_valid_i_0_4                              (cast_valid_pe_2_nw[0][4]),
    .cast_ready_o_0_4                              (cast_ready_nw_2_pe[0][4]),
    .merge_data_i_0_4                              (merge_data_pe_2_nw[0][4]),
    .merge_valid_i_0_4                             (merge_valid_pe_2_nw[0][4]),
    .merge_ready_o_0_4                             (merge_ready_nw_2_pe[0][4]),
    .gather_data_i_0_4                             (gather_data_pe_2_nw[0][4]),
    .gather_valid_i_0_4                            (gather_valid_pe_2_nw[0][4]),
    .gather_ready_o_0_4                            (gather_ready_nw_2_pe[0][4]),

    .cast_data_o_0_4                               (cast_data_nw_2_pe[0][4]),
    .cast_valid_o_0_4                              (cast_valid_nw_2_pe[0][4]),
    .cast_ready_i_0_4                              (cast_ready_pe_2_nw[0][4]),
    .merge_data_o_0_4                              (merge_data_nw_2_pe[0][4]),
    .merge_valid_o_0_4                             (merge_valid_nw_2_pe[0][4]),
    .merge_ready_i_0_4                             (merge_ready_pe_2_nw[0][4]),
    .gather_data_o_0_4                             (gather_data_nw_2_pe[0][4]),
    .gather_valid_o_0_4                            (gather_valid_nw_2_pe[0][4]),
    .gather_ready_i_0_4                            (gather_ready_pe_2_nw[0][4]),
    .cast_data_i_0_5                               (cast_data_pe_2_nw[0][5]),
    .cast_valid_i_0_5                              (cast_valid_pe_2_nw[0][5]),
    .cast_ready_o_0_5                              (cast_ready_nw_2_pe[0][5]),
    .merge_data_i_0_5                              (merge_data_pe_2_nw[0][5]),
    .merge_valid_i_0_5                             (merge_valid_pe_2_nw[0][5]),
    .merge_ready_o_0_5                             (merge_ready_nw_2_pe[0][5]),
    .gather_data_i_0_5                             (gather_data_pe_2_nw[0][5]),
    .gather_valid_i_0_5                            (gather_valid_pe_2_nw[0][5]),
    .gather_ready_o_0_5                            (gather_ready_nw_2_pe[0][5]),

    .cast_data_o_0_5                               (cast_data_nw_2_pe[0][5]),
    .cast_valid_o_0_5                              (cast_valid_nw_2_pe[0][5]),
    .cast_ready_i_0_5                              (cast_ready_pe_2_nw[0][5]),
    .merge_data_o_0_5                              (merge_data_nw_2_pe[0][5]),
    .merge_valid_o_0_5                             (merge_valid_nw_2_pe[0][5]),
    .merge_ready_i_0_5                             (merge_ready_pe_2_nw[0][5]),
    .gather_data_o_0_5                             (gather_data_nw_2_pe[0][5]),
    .gather_valid_o_0_5                            (gather_valid_nw_2_pe[0][5]),
    .gather_ready_i_0_5                            (gather_ready_pe_2_nw[0][5]),
    .cast_data_i_0_6                               (cast_data_pe_2_nw[0][6]),
    .cast_valid_i_0_6                              (cast_valid_pe_2_nw[0][6]),
    .cast_ready_o_0_6                              (cast_ready_nw_2_pe[0][6]),
    .merge_data_i_0_6                              (merge_data_pe_2_nw[0][6]),
    .merge_valid_i_0_6                             (merge_valid_pe_2_nw[0][6]),
    .merge_ready_o_0_6                             (merge_ready_nw_2_pe[0][6]),
    .gather_data_i_0_6                             (gather_data_pe_2_nw[0][6]),
    .gather_valid_i_0_6                            (gather_valid_pe_2_nw[0][6]),
    .gather_ready_o_0_6                            (gather_ready_nw_2_pe[0][6]),

    .cast_data_o_0_6                               (cast_data_nw_2_pe[0][6]),
    .cast_valid_o_0_6                              (cast_valid_nw_2_pe[0][6]),
    .cast_ready_i_0_6                              (cast_ready_pe_2_nw[0][6]),
    .merge_data_o_0_6                              (merge_data_nw_2_pe[0][6]),
    .merge_valid_o_0_6                             (merge_valid_nw_2_pe[0][6]),
    .merge_ready_i_0_6                             (merge_ready_pe_2_nw[0][6]),
    .gather_data_o_0_6                             (gather_data_nw_2_pe[0][6]),
    .gather_valid_o_0_6                            (gather_valid_nw_2_pe[0][6]),
    .gather_ready_i_0_6                            (gather_ready_pe_2_nw[0][6]),
    .cast_data_i_0_7                               (cast_data_pe_2_nw[0][7]),
    .cast_valid_i_0_7                              (cast_valid_pe_2_nw[0][7]),
    .cast_ready_o_0_7                              (cast_ready_nw_2_pe[0][7]),
    .merge_data_i_0_7                              (merge_data_pe_2_nw[0][7]),
    .merge_valid_i_0_7                             (merge_valid_pe_2_nw[0][7]),
    .merge_ready_o_0_7                             (merge_ready_nw_2_pe[0][7]),
    .gather_data_i_0_7                             (gather_data_pe_2_nw[0][7]),
    .gather_valid_i_0_7                            (gather_valid_pe_2_nw[0][7]),
    .gather_ready_o_0_7                            (gather_ready_nw_2_pe[0][7]),

    .cast_data_o_0_7                               (cast_data_nw_2_pe[0][7]),
    .cast_valid_o_0_7                              (cast_valid_nw_2_pe[0][7]),
    .cast_ready_i_0_7                              (cast_ready_pe_2_nw[0][7]),
    .merge_data_o_0_7                              (merge_data_nw_2_pe[0][7]),
    .merge_valid_o_0_7                             (merge_valid_nw_2_pe[0][7]),
    .merge_ready_i_0_7                             (merge_ready_pe_2_nw[0][7]),
    .gather_data_o_0_7                             (gather_data_nw_2_pe[0][7]),
    .gather_valid_o_0_7                            (gather_valid_nw_2_pe[0][7]),
    .gather_ready_i_0_7                            (gather_ready_pe_2_nw[0][7]),
    .cast_data_i_0_8                               (cast_data_pe_2_nw[0][8]),
    .cast_valid_i_0_8                              (cast_valid_pe_2_nw[0][8]),
    .cast_ready_o_0_8                              (cast_ready_nw_2_pe[0][8]),
    .merge_data_i_0_8                              (merge_data_pe_2_nw[0][8]),
    .merge_valid_i_0_8                             (merge_valid_pe_2_nw[0][8]),
    .merge_ready_o_0_8                             (merge_ready_nw_2_pe[0][8]),
    .gather_data_i_0_8                             (gather_data_pe_2_nw[0][8]),
    .gather_valid_i_0_8                            (gather_valid_pe_2_nw[0][8]),
    .gather_ready_o_0_8                            (gather_ready_nw_2_pe[0][8]),

    .cast_data_o_0_8                               (cast_data_nw_2_pe[0][8]),
    .cast_valid_o_0_8                              (cast_valid_nw_2_pe[0][8]),
    .cast_ready_i_0_8                              (cast_ready_pe_2_nw[0][8]),
    .merge_data_o_0_8                              (merge_data_nw_2_pe[0][8]),
    .merge_valid_o_0_8                             (merge_valid_nw_2_pe[0][8]),
    .merge_ready_i_0_8                             (merge_ready_pe_2_nw[0][8]),
    .gather_data_o_0_8                             (gather_data_nw_2_pe[0][8]),
    .gather_valid_o_0_8                            (gather_valid_nw_2_pe[0][8]),
    .gather_ready_i_0_8                            (gather_ready_pe_2_nw[0][8]),
    .cast_data_i_0_9                               (cast_data_pe_2_nw[0][9]),
    .cast_valid_i_0_9                              (cast_valid_pe_2_nw[0][9]),
    .cast_ready_o_0_9                              (cast_ready_nw_2_pe[0][9]),
    .merge_data_i_0_9                              (merge_data_pe_2_nw[0][9]),
    .merge_valid_i_0_9                             (merge_valid_pe_2_nw[0][9]),
    .merge_ready_o_0_9                             (merge_ready_nw_2_pe[0][9]),
    .gather_data_i_0_9                             (gather_data_pe_2_nw[0][9]),
    .gather_valid_i_0_9                            (gather_valid_pe_2_nw[0][9]),
    .gather_ready_o_0_9                            (gather_ready_nw_2_pe[0][9]),

    .cast_data_o_0_9                               (cast_data_nw_2_pe[0][9]),
    .cast_valid_o_0_9                              (cast_valid_nw_2_pe[0][9]),
    .cast_ready_i_0_9                              (cast_ready_pe_2_nw[0][9]),
    .merge_data_o_0_9                              (merge_data_nw_2_pe[0][9]),
    .merge_valid_o_0_9                             (merge_valid_nw_2_pe[0][9]),
    .merge_ready_i_0_9                             (merge_ready_pe_2_nw[0][9]),
    .gather_data_o_0_9                             (gather_data_nw_2_pe[0][9]),
    .gather_valid_o_0_9                            (gather_valid_nw_2_pe[0][9]),
    .gather_ready_i_0_9                            (gather_ready_pe_2_nw[0][9]),
    .cast_data_i_1_0                               (cast_data_pe_2_nw[1][0]),
    .cast_valid_i_1_0                              (cast_valid_pe_2_nw[1][0]),
    .cast_ready_o_1_0                              (cast_ready_nw_2_pe[1][0]),
    .merge_data_i_1_0                              (merge_data_pe_2_nw[1][0]),
    .merge_valid_i_1_0                             (merge_valid_pe_2_nw[1][0]),
    .merge_ready_o_1_0                             (merge_ready_nw_2_pe[1][0]),
    .gather_data_i_1_0                             (gather_data_pe_2_nw[1][0]),
    .gather_valid_i_1_0                            (gather_valid_pe_2_nw[1][0]),
    .gather_ready_o_1_0                            (gather_ready_nw_2_pe[1][0]),

    .cast_data_o_1_0                               (cast_data_nw_2_pe[1][0]),
    .cast_valid_o_1_0                              (cast_valid_nw_2_pe[1][0]),
    .cast_ready_i_1_0                              (cast_ready_pe_2_nw[1][0]),
    .merge_data_o_1_0                              (merge_data_nw_2_pe[1][0]),
    .merge_valid_o_1_0                             (merge_valid_nw_2_pe[1][0]),
    .merge_ready_i_1_0                             (merge_ready_pe_2_nw[1][0]),
    .gather_data_o_1_0                             (gather_data_nw_2_pe[1][0]),
    .gather_valid_o_1_0                            (gather_valid_nw_2_pe[1][0]),
    .gather_ready_i_1_0                            (gather_ready_pe_2_nw[1][0]),
    .cast_data_i_1_1                               (cast_data_pe_2_nw[1][1]),
    .cast_valid_i_1_1                              (cast_valid_pe_2_nw[1][1]),
    .cast_ready_o_1_1                              (cast_ready_nw_2_pe[1][1]),
    .merge_data_i_1_1                              (merge_data_pe_2_nw[1][1]),
    .merge_valid_i_1_1                             (merge_valid_pe_2_nw[1][1]),
    .merge_ready_o_1_1                             (merge_ready_nw_2_pe[1][1]),
    .gather_data_i_1_1                             (gather_data_pe_2_nw[1][1]),
    .gather_valid_i_1_1                            (gather_valid_pe_2_nw[1][1]),
    .gather_ready_o_1_1                            (gather_ready_nw_2_pe[1][1]),

    .cast_data_o_1_1                               (cast_data_nw_2_pe[1][1]),
    .cast_valid_o_1_1                              (cast_valid_nw_2_pe[1][1]),
    .cast_ready_i_1_1                              (cast_ready_pe_2_nw[1][1]),
    .merge_data_o_1_1                              (merge_data_nw_2_pe[1][1]),
    .merge_valid_o_1_1                             (merge_valid_nw_2_pe[1][1]),
    .merge_ready_i_1_1                             (merge_ready_pe_2_nw[1][1]),
    .gather_data_o_1_1                             (gather_data_nw_2_pe[1][1]),
    .gather_valid_o_1_1                            (gather_valid_nw_2_pe[1][1]),
    .gather_ready_i_1_1                            (gather_ready_pe_2_nw[1][1]),
    .cast_data_i_1_2                               (cast_data_pe_2_nw[1][2]),
    .cast_valid_i_1_2                              (cast_valid_pe_2_nw[1][2]),
    .cast_ready_o_1_2                              (cast_ready_nw_2_pe[1][2]),
    .merge_data_i_1_2                              (merge_data_pe_2_nw[1][2]),
    .merge_valid_i_1_2                             (merge_valid_pe_2_nw[1][2]),
    .merge_ready_o_1_2                             (merge_ready_nw_2_pe[1][2]),
    .gather_data_i_1_2                             (gather_data_pe_2_nw[1][2]),
    .gather_valid_i_1_2                            (gather_valid_pe_2_nw[1][2]),
    .gather_ready_o_1_2                            (gather_ready_nw_2_pe[1][2]),

    .cast_data_o_1_2                               (cast_data_nw_2_pe[1][2]),
    .cast_valid_o_1_2                              (cast_valid_nw_2_pe[1][2]),
    .cast_ready_i_1_2                              (cast_ready_pe_2_nw[1][2]),
    .merge_data_o_1_2                              (merge_data_nw_2_pe[1][2]),
    .merge_valid_o_1_2                             (merge_valid_nw_2_pe[1][2]),
    .merge_ready_i_1_2                             (merge_ready_pe_2_nw[1][2]),
    .gather_data_o_1_2                             (gather_data_nw_2_pe[1][2]),
    .gather_valid_o_1_2                            (gather_valid_nw_2_pe[1][2]),
    .gather_ready_i_1_2                            (gather_ready_pe_2_nw[1][2]),
    .cast_data_i_1_3                               (cast_data_pe_2_nw[1][3]),
    .cast_valid_i_1_3                              (cast_valid_pe_2_nw[1][3]),
    .cast_ready_o_1_3                              (cast_ready_nw_2_pe[1][3]),
    .merge_data_i_1_3                              (merge_data_pe_2_nw[1][3]),
    .merge_valid_i_1_3                             (merge_valid_pe_2_nw[1][3]),
    .merge_ready_o_1_3                             (merge_ready_nw_2_pe[1][3]),
    .gather_data_i_1_3                             (gather_data_pe_2_nw[1][3]),
    .gather_valid_i_1_3                            (gather_valid_pe_2_nw[1][3]),
    .gather_ready_o_1_3                            (gather_ready_nw_2_pe[1][3]),

    .cast_data_o_1_3                               (cast_data_nw_2_pe[1][3]),
    .cast_valid_o_1_3                              (cast_valid_nw_2_pe[1][3]),
    .cast_ready_i_1_3                              (cast_ready_pe_2_nw[1][3]),
    .merge_data_o_1_3                              (merge_data_nw_2_pe[1][3]),
    .merge_valid_o_1_3                             (merge_valid_nw_2_pe[1][3]),
    .merge_ready_i_1_3                             (merge_ready_pe_2_nw[1][3]),
    .gather_data_o_1_3                             (gather_data_nw_2_pe[1][3]),
    .gather_valid_o_1_3                            (gather_valid_nw_2_pe[1][3]),
    .gather_ready_i_1_3                            (gather_ready_pe_2_nw[1][3]),
    .cast_data_i_1_4                               (cast_data_pe_2_nw[1][4]),
    .cast_valid_i_1_4                              (cast_valid_pe_2_nw[1][4]),
    .cast_ready_o_1_4                              (cast_ready_nw_2_pe[1][4]),
    .merge_data_i_1_4                              (merge_data_pe_2_nw[1][4]),
    .merge_valid_i_1_4                             (merge_valid_pe_2_nw[1][4]),
    .merge_ready_o_1_4                             (merge_ready_nw_2_pe[1][4]),
    .gather_data_i_1_4                             (gather_data_pe_2_nw[1][4]),
    .gather_valid_i_1_4                            (gather_valid_pe_2_nw[1][4]),
    .gather_ready_o_1_4                            (gather_ready_nw_2_pe[1][4]),

    .cast_data_o_1_4                               (cast_data_nw_2_pe[1][4]),
    .cast_valid_o_1_4                              (cast_valid_nw_2_pe[1][4]),
    .cast_ready_i_1_4                              (cast_ready_pe_2_nw[1][4]),
    .merge_data_o_1_4                              (merge_data_nw_2_pe[1][4]),
    .merge_valid_o_1_4                             (merge_valid_nw_2_pe[1][4]),
    .merge_ready_i_1_4                             (merge_ready_pe_2_nw[1][4]),
    .gather_data_o_1_4                             (gather_data_nw_2_pe[1][4]),
    .gather_valid_o_1_4                            (gather_valid_nw_2_pe[1][4]),
    .gather_ready_i_1_4                            (gather_ready_pe_2_nw[1][4]),
    .cast_data_i_1_5                               (cast_data_pe_2_nw[1][5]),
    .cast_valid_i_1_5                              (cast_valid_pe_2_nw[1][5]),
    .cast_ready_o_1_5                              (cast_ready_nw_2_pe[1][5]),
    .merge_data_i_1_5                              (merge_data_pe_2_nw[1][5]),
    .merge_valid_i_1_5                             (merge_valid_pe_2_nw[1][5]),
    .merge_ready_o_1_5                             (merge_ready_nw_2_pe[1][5]),
    .gather_data_i_1_5                             (gather_data_pe_2_nw[1][5]),
    .gather_valid_i_1_5                            (gather_valid_pe_2_nw[1][5]),
    .gather_ready_o_1_5                            (gather_ready_nw_2_pe[1][5]),

    .cast_data_o_1_5                               (cast_data_nw_2_pe[1][5]),
    .cast_valid_o_1_5                              (cast_valid_nw_2_pe[1][5]),
    .cast_ready_i_1_5                              (cast_ready_pe_2_nw[1][5]),
    .merge_data_o_1_5                              (merge_data_nw_2_pe[1][5]),
    .merge_valid_o_1_5                             (merge_valid_nw_2_pe[1][5]),
    .merge_ready_i_1_5                             (merge_ready_pe_2_nw[1][5]),
    .gather_data_o_1_5                             (gather_data_nw_2_pe[1][5]),
    .gather_valid_o_1_5                            (gather_valid_nw_2_pe[1][5]),
    .gather_ready_i_1_5                            (gather_ready_pe_2_nw[1][5]),
    .cast_data_i_1_6                               (cast_data_pe_2_nw[1][6]),
    .cast_valid_i_1_6                              (cast_valid_pe_2_nw[1][6]),
    .cast_ready_o_1_6                              (cast_ready_nw_2_pe[1][6]),
    .merge_data_i_1_6                              (merge_data_pe_2_nw[1][6]),
    .merge_valid_i_1_6                             (merge_valid_pe_2_nw[1][6]),
    .merge_ready_o_1_6                             (merge_ready_nw_2_pe[1][6]),
    .gather_data_i_1_6                             (gather_data_pe_2_nw[1][6]),
    .gather_valid_i_1_6                            (gather_valid_pe_2_nw[1][6]),
    .gather_ready_o_1_6                            (gather_ready_nw_2_pe[1][6]),

    .cast_data_o_1_6                               (cast_data_nw_2_pe[1][6]),
    .cast_valid_o_1_6                              (cast_valid_nw_2_pe[1][6]),
    .cast_ready_i_1_6                              (cast_ready_pe_2_nw[1][6]),
    .merge_data_o_1_6                              (merge_data_nw_2_pe[1][6]),
    .merge_valid_o_1_6                             (merge_valid_nw_2_pe[1][6]),
    .merge_ready_i_1_6                             (merge_ready_pe_2_nw[1][6]),
    .gather_data_o_1_6                             (gather_data_nw_2_pe[1][6]),
    .gather_valid_o_1_6                            (gather_valid_nw_2_pe[1][6]),
    .gather_ready_i_1_6                            (gather_ready_pe_2_nw[1][6]),
    .cast_data_i_1_7                               (cast_data_pe_2_nw[1][7]),
    .cast_valid_i_1_7                              (cast_valid_pe_2_nw[1][7]),
    .cast_ready_o_1_7                              (cast_ready_nw_2_pe[1][7]),
    .merge_data_i_1_7                              (merge_data_pe_2_nw[1][7]),
    .merge_valid_i_1_7                             (merge_valid_pe_2_nw[1][7]),
    .merge_ready_o_1_7                             (merge_ready_nw_2_pe[1][7]),
    .gather_data_i_1_7                             (gather_data_pe_2_nw[1][7]),
    .gather_valid_i_1_7                            (gather_valid_pe_2_nw[1][7]),
    .gather_ready_o_1_7                            (gather_ready_nw_2_pe[1][7]),

    .cast_data_o_1_7                               (cast_data_nw_2_pe[1][7]),
    .cast_valid_o_1_7                              (cast_valid_nw_2_pe[1][7]),
    .cast_ready_i_1_7                              (cast_ready_pe_2_nw[1][7]),
    .merge_data_o_1_7                              (merge_data_nw_2_pe[1][7]),
    .merge_valid_o_1_7                             (merge_valid_nw_2_pe[1][7]),
    .merge_ready_i_1_7                             (merge_ready_pe_2_nw[1][7]),
    .gather_data_o_1_7                             (gather_data_nw_2_pe[1][7]),
    .gather_valid_o_1_7                            (gather_valid_nw_2_pe[1][7]),
    .gather_ready_i_1_7                            (gather_ready_pe_2_nw[1][7]),
    .cast_data_i_1_8                               (cast_data_pe_2_nw[1][8]),
    .cast_valid_i_1_8                              (cast_valid_pe_2_nw[1][8]),
    .cast_ready_o_1_8                              (cast_ready_nw_2_pe[1][8]),
    .merge_data_i_1_8                              (merge_data_pe_2_nw[1][8]),
    .merge_valid_i_1_8                             (merge_valid_pe_2_nw[1][8]),
    .merge_ready_o_1_8                             (merge_ready_nw_2_pe[1][8]),
    .gather_data_i_1_8                             (gather_data_pe_2_nw[1][8]),
    .gather_valid_i_1_8                            (gather_valid_pe_2_nw[1][8]),
    .gather_ready_o_1_8                            (gather_ready_nw_2_pe[1][8]),

    .cast_data_o_1_8                               (cast_data_nw_2_pe[1][8]),
    .cast_valid_o_1_8                              (cast_valid_nw_2_pe[1][8]),
    .cast_ready_i_1_8                              (cast_ready_pe_2_nw[1][8]),
    .merge_data_o_1_8                              (merge_data_nw_2_pe[1][8]),
    .merge_valid_o_1_8                             (merge_valid_nw_2_pe[1][8]),
    .merge_ready_i_1_8                             (merge_ready_pe_2_nw[1][8]),
    .gather_data_o_1_8                             (gather_data_nw_2_pe[1][8]),
    .gather_valid_o_1_8                            (gather_valid_nw_2_pe[1][8]),
    .gather_ready_i_1_8                            (gather_ready_pe_2_nw[1][8]),
    .cast_data_i_1_9                               (cast_data_pe_2_nw[1][9]),
    .cast_valid_i_1_9                              (cast_valid_pe_2_nw[1][9]),
    .cast_ready_o_1_9                              (cast_ready_nw_2_pe[1][9]),
    .merge_data_i_1_9                              (merge_data_pe_2_nw[1][9]),
    .merge_valid_i_1_9                             (merge_valid_pe_2_nw[1][9]),
    .merge_ready_o_1_9                             (merge_ready_nw_2_pe[1][9]),
    .gather_data_i_1_9                             (gather_data_pe_2_nw[1][9]),
    .gather_valid_i_1_9                            (gather_valid_pe_2_nw[1][9]),
    .gather_ready_o_1_9                            (gather_ready_nw_2_pe[1][9]),

    .cast_data_o_1_9                               (cast_data_nw_2_pe[1][9]),
    .cast_valid_o_1_9                              (cast_valid_nw_2_pe[1][9]),
    .cast_ready_i_1_9                              (cast_ready_pe_2_nw[1][9]),
    .merge_data_o_1_9                              (merge_data_nw_2_pe[1][9]),
    .merge_valid_o_1_9                             (merge_valid_nw_2_pe[1][9]),
    .merge_ready_i_1_9                             (merge_ready_pe_2_nw[1][9]),
    .gather_data_o_1_9                             (gather_data_nw_2_pe[1][9]),
    .gather_valid_o_1_9                            (gather_valid_nw_2_pe[1][9]),
    .gather_ready_i_1_9                            (gather_ready_pe_2_nw[1][9]),
    .cast_data_i_2_0                               (cast_data_pe_2_nw[2][0]),
    .cast_valid_i_2_0                              (cast_valid_pe_2_nw[2][0]),
    .cast_ready_o_2_0                              (cast_ready_nw_2_pe[2][0]),
    .merge_data_i_2_0                              (merge_data_pe_2_nw[2][0]),
    .merge_valid_i_2_0                             (merge_valid_pe_2_nw[2][0]),
    .merge_ready_o_2_0                             (merge_ready_nw_2_pe[2][0]),
    .gather_data_i_2_0                             (gather_data_pe_2_nw[2][0]),
    .gather_valid_i_2_0                            (gather_valid_pe_2_nw[2][0]),
    .gather_ready_o_2_0                            (gather_ready_nw_2_pe[2][0]),

    .cast_data_o_2_0                               (cast_data_nw_2_pe[2][0]),
    .cast_valid_o_2_0                              (cast_valid_nw_2_pe[2][0]),
    .cast_ready_i_2_0                              (cast_ready_pe_2_nw[2][0]),
    .merge_data_o_2_0                              (merge_data_nw_2_pe[2][0]),
    .merge_valid_o_2_0                             (merge_valid_nw_2_pe[2][0]),
    .merge_ready_i_2_0                             (merge_ready_pe_2_nw[2][0]),
    .gather_data_o_2_0                             (gather_data_nw_2_pe[2][0]),
    .gather_valid_o_2_0                            (gather_valid_nw_2_pe[2][0]),
    .gather_ready_i_2_0                            (gather_ready_pe_2_nw[2][0]),
    .cast_data_i_2_1                               (cast_data_pe_2_nw[2][1]),
    .cast_valid_i_2_1                              (cast_valid_pe_2_nw[2][1]),
    .cast_ready_o_2_1                              (cast_ready_nw_2_pe[2][1]),
    .merge_data_i_2_1                              (merge_data_pe_2_nw[2][1]),
    .merge_valid_i_2_1                             (merge_valid_pe_2_nw[2][1]),
    .merge_ready_o_2_1                             (merge_ready_nw_2_pe[2][1]),
    .gather_data_i_2_1                             (gather_data_pe_2_nw[2][1]),
    .gather_valid_i_2_1                            (gather_valid_pe_2_nw[2][1]),
    .gather_ready_o_2_1                            (gather_ready_nw_2_pe[2][1]),

    .cast_data_o_2_1                               (cast_data_nw_2_pe[2][1]),
    .cast_valid_o_2_1                              (cast_valid_nw_2_pe[2][1]),
    .cast_ready_i_2_1                              (cast_ready_pe_2_nw[2][1]),
    .merge_data_o_2_1                              (merge_data_nw_2_pe[2][1]),
    .merge_valid_o_2_1                             (merge_valid_nw_2_pe[2][1]),
    .merge_ready_i_2_1                             (merge_ready_pe_2_nw[2][1]),
    .gather_data_o_2_1                             (gather_data_nw_2_pe[2][1]),
    .gather_valid_o_2_1                            (gather_valid_nw_2_pe[2][1]),
    .gather_ready_i_2_1                            (gather_ready_pe_2_nw[2][1]),
    .cast_data_i_2_2                               (cast_data_pe_2_nw[2][2]),
    .cast_valid_i_2_2                              (cast_valid_pe_2_nw[2][2]),
    .cast_ready_o_2_2                              (cast_ready_nw_2_pe[2][2]),
    .merge_data_i_2_2                              (merge_data_pe_2_nw[2][2]),
    .merge_valid_i_2_2                             (merge_valid_pe_2_nw[2][2]),
    .merge_ready_o_2_2                             (merge_ready_nw_2_pe[2][2]),
    .gather_data_i_2_2                             (gather_data_pe_2_nw[2][2]),
    .gather_valid_i_2_2                            (gather_valid_pe_2_nw[2][2]),
    .gather_ready_o_2_2                            (gather_ready_nw_2_pe[2][2]),

    .cast_data_o_2_2                               (cast_data_nw_2_pe[2][2]),
    .cast_valid_o_2_2                              (cast_valid_nw_2_pe[2][2]),
    .cast_ready_i_2_2                              (cast_ready_pe_2_nw[2][2]),
    .merge_data_o_2_2                              (merge_data_nw_2_pe[2][2]),
    .merge_valid_o_2_2                             (merge_valid_nw_2_pe[2][2]),
    .merge_ready_i_2_2                             (merge_ready_pe_2_nw[2][2]),
    .gather_data_o_2_2                             (gather_data_nw_2_pe[2][2]),
    .gather_valid_o_2_2                            (gather_valid_nw_2_pe[2][2]),
    .gather_ready_i_2_2                            (gather_ready_pe_2_nw[2][2]),
    .cast_data_i_2_3                               (cast_data_pe_2_nw[2][3]),
    .cast_valid_i_2_3                              (cast_valid_pe_2_nw[2][3]),
    .cast_ready_o_2_3                              (cast_ready_nw_2_pe[2][3]),
    .merge_data_i_2_3                              (merge_data_pe_2_nw[2][3]),
    .merge_valid_i_2_3                             (merge_valid_pe_2_nw[2][3]),
    .merge_ready_o_2_3                             (merge_ready_nw_2_pe[2][3]),
    .gather_data_i_2_3                             (gather_data_pe_2_nw[2][3]),
    .gather_valid_i_2_3                            (gather_valid_pe_2_nw[2][3]),
    .gather_ready_o_2_3                            (gather_ready_nw_2_pe[2][3]),

    .cast_data_o_2_3                               (cast_data_nw_2_pe[2][3]),
    .cast_valid_o_2_3                              (cast_valid_nw_2_pe[2][3]),
    .cast_ready_i_2_3                              (cast_ready_pe_2_nw[2][3]),
    .merge_data_o_2_3                              (merge_data_nw_2_pe[2][3]),
    .merge_valid_o_2_3                             (merge_valid_nw_2_pe[2][3]),
    .merge_ready_i_2_3                             (merge_ready_pe_2_nw[2][3]),
    .gather_data_o_2_3                             (gather_data_nw_2_pe[2][3]),
    .gather_valid_o_2_3                            (gather_valid_nw_2_pe[2][3]),
    .gather_ready_i_2_3                            (gather_ready_pe_2_nw[2][3]),
    .cast_data_i_2_4                               (cast_data_pe_2_nw[2][4]),
    .cast_valid_i_2_4                              (cast_valid_pe_2_nw[2][4]),
    .cast_ready_o_2_4                              (cast_ready_nw_2_pe[2][4]),
    .merge_data_i_2_4                              (merge_data_pe_2_nw[2][4]),
    .merge_valid_i_2_4                             (merge_valid_pe_2_nw[2][4]),
    .merge_ready_o_2_4                             (merge_ready_nw_2_pe[2][4]),
    .gather_data_i_2_4                             (gather_data_pe_2_nw[2][4]),
    .gather_valid_i_2_4                            (gather_valid_pe_2_nw[2][4]),
    .gather_ready_o_2_4                            (gather_ready_nw_2_pe[2][4]),

    .cast_data_o_2_4                               (cast_data_nw_2_pe[2][4]),
    .cast_valid_o_2_4                              (cast_valid_nw_2_pe[2][4]),
    .cast_ready_i_2_4                              (cast_ready_pe_2_nw[2][4]),
    .merge_data_o_2_4                              (merge_data_nw_2_pe[2][4]),
    .merge_valid_o_2_4                             (merge_valid_nw_2_pe[2][4]),
    .merge_ready_i_2_4                             (merge_ready_pe_2_nw[2][4]),
    .gather_data_o_2_4                             (gather_data_nw_2_pe[2][4]),
    .gather_valid_o_2_4                            (gather_valid_nw_2_pe[2][4]),
    .gather_ready_i_2_4                            (gather_ready_pe_2_nw[2][4]),
    .cast_data_i_2_5                               (cast_data_pe_2_nw[2][5]),
    .cast_valid_i_2_5                              (cast_valid_pe_2_nw[2][5]),
    .cast_ready_o_2_5                              (cast_ready_nw_2_pe[2][5]),
    .merge_data_i_2_5                              (merge_data_pe_2_nw[2][5]),
    .merge_valid_i_2_5                             (merge_valid_pe_2_nw[2][5]),
    .merge_ready_o_2_5                             (merge_ready_nw_2_pe[2][5]),
    .gather_data_i_2_5                             (gather_data_pe_2_nw[2][5]),
    .gather_valid_i_2_5                            (gather_valid_pe_2_nw[2][5]),
    .gather_ready_o_2_5                            (gather_ready_nw_2_pe[2][5]),

    .cast_data_o_2_5                               (cast_data_nw_2_pe[2][5]),
    .cast_valid_o_2_5                              (cast_valid_nw_2_pe[2][5]),
    .cast_ready_i_2_5                              (cast_ready_pe_2_nw[2][5]),
    .merge_data_o_2_5                              (merge_data_nw_2_pe[2][5]),
    .merge_valid_o_2_5                             (merge_valid_nw_2_pe[2][5]),
    .merge_ready_i_2_5                             (merge_ready_pe_2_nw[2][5]),
    .gather_data_o_2_5                             (gather_data_nw_2_pe[2][5]),
    .gather_valid_o_2_5                            (gather_valid_nw_2_pe[2][5]),
    .gather_ready_i_2_5                            (gather_ready_pe_2_nw[2][5]),
    .cast_data_i_2_6                               (cast_data_pe_2_nw[2][6]),
    .cast_valid_i_2_6                              (cast_valid_pe_2_nw[2][6]),
    .cast_ready_o_2_6                              (cast_ready_nw_2_pe[2][6]),
    .merge_data_i_2_6                              (merge_data_pe_2_nw[2][6]),
    .merge_valid_i_2_6                             (merge_valid_pe_2_nw[2][6]),
    .merge_ready_o_2_6                             (merge_ready_nw_2_pe[2][6]),
    .gather_data_i_2_6                             (gather_data_pe_2_nw[2][6]),
    .gather_valid_i_2_6                            (gather_valid_pe_2_nw[2][6]),
    .gather_ready_o_2_6                            (gather_ready_nw_2_pe[2][6]),

    .cast_data_o_2_6                               (cast_data_nw_2_pe[2][6]),
    .cast_valid_o_2_6                              (cast_valid_nw_2_pe[2][6]),
    .cast_ready_i_2_6                              (cast_ready_pe_2_nw[2][6]),
    .merge_data_o_2_6                              (merge_data_nw_2_pe[2][6]),
    .merge_valid_o_2_6                             (merge_valid_nw_2_pe[2][6]),
    .merge_ready_i_2_6                             (merge_ready_pe_2_nw[2][6]),
    .gather_data_o_2_6                             (gather_data_nw_2_pe[2][6]),
    .gather_valid_o_2_6                            (gather_valid_nw_2_pe[2][6]),
    .gather_ready_i_2_6                            (gather_ready_pe_2_nw[2][6]),
    .cast_data_i_2_7                               (cast_data_pe_2_nw[2][7]),
    .cast_valid_i_2_7                              (cast_valid_pe_2_nw[2][7]),
    .cast_ready_o_2_7                              (cast_ready_nw_2_pe[2][7]),
    .merge_data_i_2_7                              (merge_data_pe_2_nw[2][7]),
    .merge_valid_i_2_7                             (merge_valid_pe_2_nw[2][7]),
    .merge_ready_o_2_7                             (merge_ready_nw_2_pe[2][7]),
    .gather_data_i_2_7                             (gather_data_pe_2_nw[2][7]),
    .gather_valid_i_2_7                            (gather_valid_pe_2_nw[2][7]),
    .gather_ready_o_2_7                            (gather_ready_nw_2_pe[2][7]),

    .cast_data_o_2_7                               (cast_data_nw_2_pe[2][7]),
    .cast_valid_o_2_7                              (cast_valid_nw_2_pe[2][7]),
    .cast_ready_i_2_7                              (cast_ready_pe_2_nw[2][7]),
    .merge_data_o_2_7                              (merge_data_nw_2_pe[2][7]),
    .merge_valid_o_2_7                             (merge_valid_nw_2_pe[2][7]),
    .merge_ready_i_2_7                             (merge_ready_pe_2_nw[2][7]),
    .gather_data_o_2_7                             (gather_data_nw_2_pe[2][7]),
    .gather_valid_o_2_7                            (gather_valid_nw_2_pe[2][7]),
    .gather_ready_i_2_7                            (gather_ready_pe_2_nw[2][7]),
    .cast_data_i_2_8                               (cast_data_pe_2_nw[2][8]),
    .cast_valid_i_2_8                              (cast_valid_pe_2_nw[2][8]),
    .cast_ready_o_2_8                              (cast_ready_nw_2_pe[2][8]),
    .merge_data_i_2_8                              (merge_data_pe_2_nw[2][8]),
    .merge_valid_i_2_8                             (merge_valid_pe_2_nw[2][8]),
    .merge_ready_o_2_8                             (merge_ready_nw_2_pe[2][8]),
    .gather_data_i_2_8                             (gather_data_pe_2_nw[2][8]),
    .gather_valid_i_2_8                            (gather_valid_pe_2_nw[2][8]),
    .gather_ready_o_2_8                            (gather_ready_nw_2_pe[2][8]),

    .cast_data_o_2_8                               (cast_data_nw_2_pe[2][8]),
    .cast_valid_o_2_8                              (cast_valid_nw_2_pe[2][8]),
    .cast_ready_i_2_8                              (cast_ready_pe_2_nw[2][8]),
    .merge_data_o_2_8                              (merge_data_nw_2_pe[2][8]),
    .merge_valid_o_2_8                             (merge_valid_nw_2_pe[2][8]),
    .merge_ready_i_2_8                             (merge_ready_pe_2_nw[2][8]),
    .gather_data_o_2_8                             (gather_data_nw_2_pe[2][8]),
    .gather_valid_o_2_8                            (gather_valid_nw_2_pe[2][8]),
    .gather_ready_i_2_8                            (gather_ready_pe_2_nw[2][8]),
    .cast_data_i_2_9                               (cast_data_pe_2_nw[2][9]),
    .cast_valid_i_2_9                              (cast_valid_pe_2_nw[2][9]),
    .cast_ready_o_2_9                              (cast_ready_nw_2_pe[2][9]),
    .merge_data_i_2_9                              (merge_data_pe_2_nw[2][9]),
    .merge_valid_i_2_9                             (merge_valid_pe_2_nw[2][9]),
    .merge_ready_o_2_9                             (merge_ready_nw_2_pe[2][9]),
    .gather_data_i_2_9                             (gather_data_pe_2_nw[2][9]),
    .gather_valid_i_2_9                            (gather_valid_pe_2_nw[2][9]),
    .gather_ready_o_2_9                            (gather_ready_nw_2_pe[2][9]),

    .cast_data_o_2_9                               (cast_data_nw_2_pe[2][9]),
    .cast_valid_o_2_9                              (cast_valid_nw_2_pe[2][9]),
    .cast_ready_i_2_9                              (cast_ready_pe_2_nw[2][9]),
    .merge_data_o_2_9                              (merge_data_nw_2_pe[2][9]),
    .merge_valid_o_2_9                             (merge_valid_nw_2_pe[2][9]),
    .merge_ready_i_2_9                             (merge_ready_pe_2_nw[2][9]),
    .gather_data_o_2_9                             (gather_data_nw_2_pe[2][9]),
    .gather_valid_o_2_9                            (gather_valid_nw_2_pe[2][9]),
    .gather_ready_i_2_9                            (gather_ready_pe_2_nw[2][9]),
    .cast_data_i_3_0                               (cast_data_pe_2_nw[3][0]),
    .cast_valid_i_3_0                              (cast_valid_pe_2_nw[3][0]),
    .cast_ready_o_3_0                              (cast_ready_nw_2_pe[3][0]),
    .merge_data_i_3_0                              (merge_data_pe_2_nw[3][0]),
    .merge_valid_i_3_0                             (merge_valid_pe_2_nw[3][0]),
    .merge_ready_o_3_0                             (merge_ready_nw_2_pe[3][0]),
    .gather_data_i_3_0                             (gather_data_pe_2_nw[3][0]),
    .gather_valid_i_3_0                            (gather_valid_pe_2_nw[3][0]),
    .gather_ready_o_3_0                            (gather_ready_nw_2_pe[3][0]),

    .cast_data_o_3_0                               (cast_data_nw_2_pe[3][0]),
    .cast_valid_o_3_0                              (cast_valid_nw_2_pe[3][0]),
    .cast_ready_i_3_0                              (cast_ready_pe_2_nw[3][0]),
    .merge_data_o_3_0                              (merge_data_nw_2_pe[3][0]),
    .merge_valid_o_3_0                             (merge_valid_nw_2_pe[3][0]),
    .merge_ready_i_3_0                             (merge_ready_pe_2_nw[3][0]),
    .gather_data_o_3_0                             (gather_data_nw_2_pe[3][0]),
    .gather_valid_o_3_0                            (gather_valid_nw_2_pe[3][0]),
    .gather_ready_i_3_0                            (gather_ready_pe_2_nw[3][0]),
    .cast_data_i_3_1                               (cast_data_pe_2_nw[3][1]),
    .cast_valid_i_3_1                              (cast_valid_pe_2_nw[3][1]),
    .cast_ready_o_3_1                              (cast_ready_nw_2_pe[3][1]),
    .merge_data_i_3_1                              (merge_data_pe_2_nw[3][1]),
    .merge_valid_i_3_1                             (merge_valid_pe_2_nw[3][1]),
    .merge_ready_o_3_1                             (merge_ready_nw_2_pe[3][1]),
    .gather_data_i_3_1                             (gather_data_pe_2_nw[3][1]),
    .gather_valid_i_3_1                            (gather_valid_pe_2_nw[3][1]),
    .gather_ready_o_3_1                            (gather_ready_nw_2_pe[3][1]),

    .cast_data_o_3_1                               (cast_data_nw_2_pe[3][1]),
    .cast_valid_o_3_1                              (cast_valid_nw_2_pe[3][1]),
    .cast_ready_i_3_1                              (cast_ready_pe_2_nw[3][1]),
    .merge_data_o_3_1                              (merge_data_nw_2_pe[3][1]),
    .merge_valid_o_3_1                             (merge_valid_nw_2_pe[3][1]),
    .merge_ready_i_3_1                             (merge_ready_pe_2_nw[3][1]),
    .gather_data_o_3_1                             (gather_data_nw_2_pe[3][1]),
    .gather_valid_o_3_1                            (gather_valid_nw_2_pe[3][1]),
    .gather_ready_i_3_1                            (gather_ready_pe_2_nw[3][1]),
    .cast_data_i_3_2                               (cast_data_pe_2_nw[3][2]),
    .cast_valid_i_3_2                              (cast_valid_pe_2_nw[3][2]),
    .cast_ready_o_3_2                              (cast_ready_nw_2_pe[3][2]),
    .merge_data_i_3_2                              (merge_data_pe_2_nw[3][2]),
    .merge_valid_i_3_2                             (merge_valid_pe_2_nw[3][2]),
    .merge_ready_o_3_2                             (merge_ready_nw_2_pe[3][2]),
    .gather_data_i_3_2                             (gather_data_pe_2_nw[3][2]),
    .gather_valid_i_3_2                            (gather_valid_pe_2_nw[3][2]),
    .gather_ready_o_3_2                            (gather_ready_nw_2_pe[3][2]),

    .cast_data_o_3_2                               (cast_data_nw_2_pe[3][2]),
    .cast_valid_o_3_2                              (cast_valid_nw_2_pe[3][2]),
    .cast_ready_i_3_2                              (cast_ready_pe_2_nw[3][2]),
    .merge_data_o_3_2                              (merge_data_nw_2_pe[3][2]),
    .merge_valid_o_3_2                             (merge_valid_nw_2_pe[3][2]),
    .merge_ready_i_3_2                             (merge_ready_pe_2_nw[3][2]),
    .gather_data_o_3_2                             (gather_data_nw_2_pe[3][2]),
    .gather_valid_o_3_2                            (gather_valid_nw_2_pe[3][2]),
    .gather_ready_i_3_2                            (gather_ready_pe_2_nw[3][2]),
    .cast_data_i_3_3                               (cast_data_pe_2_nw[3][3]),
    .cast_valid_i_3_3                              (cast_valid_pe_2_nw[3][3]),
    .cast_ready_o_3_3                              (cast_ready_nw_2_pe[3][3]),
    .merge_data_i_3_3                              (merge_data_pe_2_nw[3][3]),
    .merge_valid_i_3_3                             (merge_valid_pe_2_nw[3][3]),
    .merge_ready_o_3_3                             (merge_ready_nw_2_pe[3][3]),
    .gather_data_i_3_3                             (gather_data_pe_2_nw[3][3]),
    .gather_valid_i_3_3                            (gather_valid_pe_2_nw[3][3]),
    .gather_ready_o_3_3                            (gather_ready_nw_2_pe[3][3]),

    .cast_data_o_3_3                               (cast_data_nw_2_pe[3][3]),
    .cast_valid_o_3_3                              (cast_valid_nw_2_pe[3][3]),
    .cast_ready_i_3_3                              (cast_ready_pe_2_nw[3][3]),
    .merge_data_o_3_3                              (merge_data_nw_2_pe[3][3]),
    .merge_valid_o_3_3                             (merge_valid_nw_2_pe[3][3]),
    .merge_ready_i_3_3                             (merge_ready_pe_2_nw[3][3]),
    .gather_data_o_3_3                             (gather_data_nw_2_pe[3][3]),
    .gather_valid_o_3_3                            (gather_valid_nw_2_pe[3][3]),
    .gather_ready_i_3_3                            (gather_ready_pe_2_nw[3][3]),
    .cast_data_i_3_4                               (cast_data_pe_2_nw[3][4]),
    .cast_valid_i_3_4                              (cast_valid_pe_2_nw[3][4]),
    .cast_ready_o_3_4                              (cast_ready_nw_2_pe[3][4]),
    .merge_data_i_3_4                              (merge_data_pe_2_nw[3][4]),
    .merge_valid_i_3_4                             (merge_valid_pe_2_nw[3][4]),
    .merge_ready_o_3_4                             (merge_ready_nw_2_pe[3][4]),
    .gather_data_i_3_4                             (gather_data_pe_2_nw[3][4]),
    .gather_valid_i_3_4                            (gather_valid_pe_2_nw[3][4]),
    .gather_ready_o_3_4                            (gather_ready_nw_2_pe[3][4]),

    .cast_data_o_3_4                               (cast_data_nw_2_pe[3][4]),
    .cast_valid_o_3_4                              (cast_valid_nw_2_pe[3][4]),
    .cast_ready_i_3_4                              (cast_ready_pe_2_nw[3][4]),
    .merge_data_o_3_4                              (merge_data_nw_2_pe[3][4]),
    .merge_valid_o_3_4                             (merge_valid_nw_2_pe[3][4]),
    .merge_ready_i_3_4                             (merge_ready_pe_2_nw[3][4]),
    .gather_data_o_3_4                             (gather_data_nw_2_pe[3][4]),
    .gather_valid_o_3_4                            (gather_valid_nw_2_pe[3][4]),
    .gather_ready_i_3_4                            (gather_ready_pe_2_nw[3][4]),
    .cast_data_i_3_5                               (cast_data_pe_2_nw[3][5]),
    .cast_valid_i_3_5                              (cast_valid_pe_2_nw[3][5]),
    .cast_ready_o_3_5                              (cast_ready_nw_2_pe[3][5]),
    .merge_data_i_3_5                              (merge_data_pe_2_nw[3][5]),
    .merge_valid_i_3_5                             (merge_valid_pe_2_nw[3][5]),
    .merge_ready_o_3_5                             (merge_ready_nw_2_pe[3][5]),
    .gather_data_i_3_5                             (gather_data_pe_2_nw[3][5]),
    .gather_valid_i_3_5                            (gather_valid_pe_2_nw[3][5]),
    .gather_ready_o_3_5                            (gather_ready_nw_2_pe[3][5]),

    .cast_data_o_3_5                               (cast_data_nw_2_pe[3][5]),
    .cast_valid_o_3_5                              (cast_valid_nw_2_pe[3][5]),
    .cast_ready_i_3_5                              (cast_ready_pe_2_nw[3][5]),
    .merge_data_o_3_5                              (merge_data_nw_2_pe[3][5]),
    .merge_valid_o_3_5                             (merge_valid_nw_2_pe[3][5]),
    .merge_ready_i_3_5                             (merge_ready_pe_2_nw[3][5]),
    .gather_data_o_3_5                             (gather_data_nw_2_pe[3][5]),
    .gather_valid_o_3_5                            (gather_valid_nw_2_pe[3][5]),
    .gather_ready_i_3_5                            (gather_ready_pe_2_nw[3][5]),
    .cast_data_i_3_6                               (cast_data_pe_2_nw[3][6]),
    .cast_valid_i_3_6                              (cast_valid_pe_2_nw[3][6]),
    .cast_ready_o_3_6                              (cast_ready_nw_2_pe[3][6]),
    .merge_data_i_3_6                              (merge_data_pe_2_nw[3][6]),
    .merge_valid_i_3_6                             (merge_valid_pe_2_nw[3][6]),
    .merge_ready_o_3_6                             (merge_ready_nw_2_pe[3][6]),
    .gather_data_i_3_6                             (gather_data_pe_2_nw[3][6]),
    .gather_valid_i_3_6                            (gather_valid_pe_2_nw[3][6]),
    .gather_ready_o_3_6                            (gather_ready_nw_2_pe[3][6]),

    .cast_data_o_3_6                               (cast_data_nw_2_pe[3][6]),
    .cast_valid_o_3_6                              (cast_valid_nw_2_pe[3][6]),
    .cast_ready_i_3_6                              (cast_ready_pe_2_nw[3][6]),
    .merge_data_o_3_6                              (merge_data_nw_2_pe[3][6]),
    .merge_valid_o_3_6                             (merge_valid_nw_2_pe[3][6]),
    .merge_ready_i_3_6                             (merge_ready_pe_2_nw[3][6]),
    .gather_data_o_3_6                             (gather_data_nw_2_pe[3][6]),
    .gather_valid_o_3_6                            (gather_valid_nw_2_pe[3][6]),
    .gather_ready_i_3_6                            (gather_ready_pe_2_nw[3][6]),
    .cast_data_i_3_7                               (cast_data_pe_2_nw[3][7]),
    .cast_valid_i_3_7                              (cast_valid_pe_2_nw[3][7]),
    .cast_ready_o_3_7                              (cast_ready_nw_2_pe[3][7]),
    .merge_data_i_3_7                              (merge_data_pe_2_nw[3][7]),
    .merge_valid_i_3_7                             (merge_valid_pe_2_nw[3][7]),
    .merge_ready_o_3_7                             (merge_ready_nw_2_pe[3][7]),
    .gather_data_i_3_7                             (gather_data_pe_2_nw[3][7]),
    .gather_valid_i_3_7                            (gather_valid_pe_2_nw[3][7]),
    .gather_ready_o_3_7                            (gather_ready_nw_2_pe[3][7]),

    .cast_data_o_3_7                               (cast_data_nw_2_pe[3][7]),
    .cast_valid_o_3_7                              (cast_valid_nw_2_pe[3][7]),
    .cast_ready_i_3_7                              (cast_ready_pe_2_nw[3][7]),
    .merge_data_o_3_7                              (merge_data_nw_2_pe[3][7]),
    .merge_valid_o_3_7                             (merge_valid_nw_2_pe[3][7]),
    .merge_ready_i_3_7                             (merge_ready_pe_2_nw[3][7]),
    .gather_data_o_3_7                             (gather_data_nw_2_pe[3][7]),
    .gather_valid_o_3_7                            (gather_valid_nw_2_pe[3][7]),
    .gather_ready_i_3_7                            (gather_ready_pe_2_nw[3][7]),
    .cast_data_i_3_8                               (cast_data_pe_2_nw[3][8]),
    .cast_valid_i_3_8                              (cast_valid_pe_2_nw[3][8]),
    .cast_ready_o_3_8                              (cast_ready_nw_2_pe[3][8]),
    .merge_data_i_3_8                              (merge_data_pe_2_nw[3][8]),
    .merge_valid_i_3_8                             (merge_valid_pe_2_nw[3][8]),
    .merge_ready_o_3_8                             (merge_ready_nw_2_pe[3][8]),
    .gather_data_i_3_8                             (gather_data_pe_2_nw[3][8]),
    .gather_valid_i_3_8                            (gather_valid_pe_2_nw[3][8]),
    .gather_ready_o_3_8                            (gather_ready_nw_2_pe[3][8]),

    .cast_data_o_3_8                               (cast_data_nw_2_pe[3][8]),
    .cast_valid_o_3_8                              (cast_valid_nw_2_pe[3][8]),
    .cast_ready_i_3_8                              (cast_ready_pe_2_nw[3][8]),
    .merge_data_o_3_8                              (merge_data_nw_2_pe[3][8]),
    .merge_valid_o_3_8                             (merge_valid_nw_2_pe[3][8]),
    .merge_ready_i_3_8                             (merge_ready_pe_2_nw[3][8]),
    .gather_data_o_3_8                             (gather_data_nw_2_pe[3][8]),
    .gather_valid_o_3_8                            (gather_valid_nw_2_pe[3][8]),
    .gather_ready_i_3_8                            (gather_ready_pe_2_nw[3][8]),
    .cast_data_i_3_9                               (cast_data_pe_2_nw[3][9]),
    .cast_valid_i_3_9                              (cast_valid_pe_2_nw[3][9]),
    .cast_ready_o_3_9                              (cast_ready_nw_2_pe[3][9]),
    .merge_data_i_3_9                              (merge_data_pe_2_nw[3][9]),
    .merge_valid_i_3_9                             (merge_valid_pe_2_nw[3][9]),
    .merge_ready_o_3_9                             (merge_ready_nw_2_pe[3][9]),
    .gather_data_i_3_9                             (gather_data_pe_2_nw[3][9]),
    .gather_valid_i_3_9                            (gather_valid_pe_2_nw[3][9]),
    .gather_ready_o_3_9                            (gather_ready_nw_2_pe[3][9]),

    .cast_data_o_3_9                               (cast_data_nw_2_pe[3][9]),
    .cast_valid_o_3_9                              (cast_valid_nw_2_pe[3][9]),
    .cast_ready_i_3_9                              (cast_ready_pe_2_nw[3][9]),
    .merge_data_o_3_9                              (merge_data_nw_2_pe[3][9]),
    .merge_valid_o_3_9                             (merge_valid_nw_2_pe[3][9]),
    .merge_ready_i_3_9                             (merge_ready_pe_2_nw[3][9]),
    .gather_data_o_3_9                             (gather_data_nw_2_pe[3][9]),
    .gather_valid_o_3_9                            (gather_valid_nw_2_pe[3][9]),
    .gather_ready_i_3_9                            (gather_ready_pe_2_nw[3][9]),
    .cast_data_i_4_0                               (cast_data_pe_2_nw[4][0]),
    .cast_valid_i_4_0                              (cast_valid_pe_2_nw[4][0]),
    .cast_ready_o_4_0                              (cast_ready_nw_2_pe[4][0]),
    .merge_data_i_4_0                              (merge_data_pe_2_nw[4][0]),
    .merge_valid_i_4_0                             (merge_valid_pe_2_nw[4][0]),
    .merge_ready_o_4_0                             (merge_ready_nw_2_pe[4][0]),
    .gather_data_i_4_0                             (gather_data_pe_2_nw[4][0]),
    .gather_valid_i_4_0                            (gather_valid_pe_2_nw[4][0]),
    .gather_ready_o_4_0                            (gather_ready_nw_2_pe[4][0]),

    .cast_data_o_4_0                               (cast_data_nw_2_pe[4][0]),
    .cast_valid_o_4_0                              (cast_valid_nw_2_pe[4][0]),
    .cast_ready_i_4_0                              (cast_ready_pe_2_nw[4][0]),
    .merge_data_o_4_0                              (merge_data_nw_2_pe[4][0]),
    .merge_valid_o_4_0                             (merge_valid_nw_2_pe[4][0]),
    .merge_ready_i_4_0                             (merge_ready_pe_2_nw[4][0]),
    .gather_data_o_4_0                             (gather_data_nw_2_pe[4][0]),
    .gather_valid_o_4_0                            (gather_valid_nw_2_pe[4][0]),
    .gather_ready_i_4_0                            (gather_ready_pe_2_nw[4][0]),
    .cast_data_i_4_1                               (cast_data_pe_2_nw[4][1]),
    .cast_valid_i_4_1                              (cast_valid_pe_2_nw[4][1]),
    .cast_ready_o_4_1                              (cast_ready_nw_2_pe[4][1]),
    .merge_data_i_4_1                              (merge_data_pe_2_nw[4][1]),
    .merge_valid_i_4_1                             (merge_valid_pe_2_nw[4][1]),
    .merge_ready_o_4_1                             (merge_ready_nw_2_pe[4][1]),
    .gather_data_i_4_1                             (gather_data_pe_2_nw[4][1]),
    .gather_valid_i_4_1                            (gather_valid_pe_2_nw[4][1]),
    .gather_ready_o_4_1                            (gather_ready_nw_2_pe[4][1]),

    .cast_data_o_4_1                               (cast_data_nw_2_pe[4][1]),
    .cast_valid_o_4_1                              (cast_valid_nw_2_pe[4][1]),
    .cast_ready_i_4_1                              (cast_ready_pe_2_nw[4][1]),
    .merge_data_o_4_1                              (merge_data_nw_2_pe[4][1]),
    .merge_valid_o_4_1                             (merge_valid_nw_2_pe[4][1]),
    .merge_ready_i_4_1                             (merge_ready_pe_2_nw[4][1]),
    .gather_data_o_4_1                             (gather_data_nw_2_pe[4][1]),
    .gather_valid_o_4_1                            (gather_valid_nw_2_pe[4][1]),
    .gather_ready_i_4_1                            (gather_ready_pe_2_nw[4][1]),
    .cast_data_i_4_2                               (cast_data_pe_2_nw[4][2]),
    .cast_valid_i_4_2                              (cast_valid_pe_2_nw[4][2]),
    .cast_ready_o_4_2                              (cast_ready_nw_2_pe[4][2]),
    .merge_data_i_4_2                              (merge_data_pe_2_nw[4][2]),
    .merge_valid_i_4_2                             (merge_valid_pe_2_nw[4][2]),
    .merge_ready_o_4_2                             (merge_ready_nw_2_pe[4][2]),
    .gather_data_i_4_2                             (gather_data_pe_2_nw[4][2]),
    .gather_valid_i_4_2                            (gather_valid_pe_2_nw[4][2]),
    .gather_ready_o_4_2                            (gather_ready_nw_2_pe[4][2]),

    .cast_data_o_4_2                               (cast_data_nw_2_pe[4][2]),
    .cast_valid_o_4_2                              (cast_valid_nw_2_pe[4][2]),
    .cast_ready_i_4_2                              (cast_ready_pe_2_nw[4][2]),
    .merge_data_o_4_2                              (merge_data_nw_2_pe[4][2]),
    .merge_valid_o_4_2                             (merge_valid_nw_2_pe[4][2]),
    .merge_ready_i_4_2                             (merge_ready_pe_2_nw[4][2]),
    .gather_data_o_4_2                             (gather_data_nw_2_pe[4][2]),
    .gather_valid_o_4_2                            (gather_valid_nw_2_pe[4][2]),
    .gather_ready_i_4_2                            (gather_ready_pe_2_nw[4][2]),
    .cast_data_i_4_3                               (cast_data_pe_2_nw[4][3]),
    .cast_valid_i_4_3                              (cast_valid_pe_2_nw[4][3]),
    .cast_ready_o_4_3                              (cast_ready_nw_2_pe[4][3]),
    .merge_data_i_4_3                              (merge_data_pe_2_nw[4][3]),
    .merge_valid_i_4_3                             (merge_valid_pe_2_nw[4][3]),
    .merge_ready_o_4_3                             (merge_ready_nw_2_pe[4][3]),
    .gather_data_i_4_3                             (gather_data_pe_2_nw[4][3]),
    .gather_valid_i_4_3                            (gather_valid_pe_2_nw[4][3]),
    .gather_ready_o_4_3                            (gather_ready_nw_2_pe[4][3]),

    .cast_data_o_4_3                               (cast_data_nw_2_pe[4][3]),
    .cast_valid_o_4_3                              (cast_valid_nw_2_pe[4][3]),
    .cast_ready_i_4_3                              (cast_ready_pe_2_nw[4][3]),
    .merge_data_o_4_3                              (merge_data_nw_2_pe[4][3]),
    .merge_valid_o_4_3                             (merge_valid_nw_2_pe[4][3]),
    .merge_ready_i_4_3                             (merge_ready_pe_2_nw[4][3]),
    .gather_data_o_4_3                             (gather_data_nw_2_pe[4][3]),
    .gather_valid_o_4_3                            (gather_valid_nw_2_pe[4][3]),
    .gather_ready_i_4_3                            (gather_ready_pe_2_nw[4][3]),
    .cast_data_i_4_4                               (cast_data_pe_2_nw[4][4]),
    .cast_valid_i_4_4                              (cast_valid_pe_2_nw[4][4]),
    .cast_ready_o_4_4                              (cast_ready_nw_2_pe[4][4]),
    .merge_data_i_4_4                              (merge_data_pe_2_nw[4][4]),
    .merge_valid_i_4_4                             (merge_valid_pe_2_nw[4][4]),
    .merge_ready_o_4_4                             (merge_ready_nw_2_pe[4][4]),
    .gather_data_i_4_4                             (gather_data_pe_2_nw[4][4]),
    .gather_valid_i_4_4                            (gather_valid_pe_2_nw[4][4]),
    .gather_ready_o_4_4                            (gather_ready_nw_2_pe[4][4]),

    .cast_data_o_4_4                               (cast_data_nw_2_pe[4][4]),
    .cast_valid_o_4_4                              (cast_valid_nw_2_pe[4][4]),
    .cast_ready_i_4_4                              (cast_ready_pe_2_nw[4][4]),
    .merge_data_o_4_4                              (merge_data_nw_2_pe[4][4]),
    .merge_valid_o_4_4                             (merge_valid_nw_2_pe[4][4]),
    .merge_ready_i_4_4                             (merge_ready_pe_2_nw[4][4]),
    .gather_data_o_4_4                             (gather_data_nw_2_pe[4][4]),
    .gather_valid_o_4_4                            (gather_valid_nw_2_pe[4][4]),
    .gather_ready_i_4_4                            (gather_ready_pe_2_nw[4][4]),
    .cast_data_i_4_5                               (cast_data_pe_2_nw[4][5]),
    .cast_valid_i_4_5                              (cast_valid_pe_2_nw[4][5]),
    .cast_ready_o_4_5                              (cast_ready_nw_2_pe[4][5]),
    .merge_data_i_4_5                              (merge_data_pe_2_nw[4][5]),
    .merge_valid_i_4_5                             (merge_valid_pe_2_nw[4][5]),
    .merge_ready_o_4_5                             (merge_ready_nw_2_pe[4][5]),
    .gather_data_i_4_5                             (gather_data_pe_2_nw[4][5]),
    .gather_valid_i_4_5                            (gather_valid_pe_2_nw[4][5]),
    .gather_ready_o_4_5                            (gather_ready_nw_2_pe[4][5]),

    .cast_data_o_4_5                               (cast_data_nw_2_pe[4][5]),
    .cast_valid_o_4_5                              (cast_valid_nw_2_pe[4][5]),
    .cast_ready_i_4_5                              (cast_ready_pe_2_nw[4][5]),
    .merge_data_o_4_5                              (merge_data_nw_2_pe[4][5]),
    .merge_valid_o_4_5                             (merge_valid_nw_2_pe[4][5]),
    .merge_ready_i_4_5                             (merge_ready_pe_2_nw[4][5]),
    .gather_data_o_4_5                             (gather_data_nw_2_pe[4][5]),
    .gather_valid_o_4_5                            (gather_valid_nw_2_pe[4][5]),
    .gather_ready_i_4_5                            (gather_ready_pe_2_nw[4][5]),
    .cast_data_i_4_6                               (cast_data_pe_2_nw[4][6]),
    .cast_valid_i_4_6                              (cast_valid_pe_2_nw[4][6]),
    .cast_ready_o_4_6                              (cast_ready_nw_2_pe[4][6]),
    .merge_data_i_4_6                              (merge_data_pe_2_nw[4][6]),
    .merge_valid_i_4_6                             (merge_valid_pe_2_nw[4][6]),
    .merge_ready_o_4_6                             (merge_ready_nw_2_pe[4][6]),
    .gather_data_i_4_6                             (gather_data_pe_2_nw[4][6]),
    .gather_valid_i_4_6                            (gather_valid_pe_2_nw[4][6]),
    .gather_ready_o_4_6                            (gather_ready_nw_2_pe[4][6]),

    .cast_data_o_4_6                               (cast_data_nw_2_pe[4][6]),
    .cast_valid_o_4_6                              (cast_valid_nw_2_pe[4][6]),
    .cast_ready_i_4_6                              (cast_ready_pe_2_nw[4][6]),
    .merge_data_o_4_6                              (merge_data_nw_2_pe[4][6]),
    .merge_valid_o_4_6                             (merge_valid_nw_2_pe[4][6]),
    .merge_ready_i_4_6                             (merge_ready_pe_2_nw[4][6]),
    .gather_data_o_4_6                             (gather_data_nw_2_pe[4][6]),
    .gather_valid_o_4_6                            (gather_valid_nw_2_pe[4][6]),
    .gather_ready_i_4_6                            (gather_ready_pe_2_nw[4][6]),
    .cast_data_i_4_7                               (cast_data_pe_2_nw[4][7]),
    .cast_valid_i_4_7                              (cast_valid_pe_2_nw[4][7]),
    .cast_ready_o_4_7                              (cast_ready_nw_2_pe[4][7]),
    .merge_data_i_4_7                              (merge_data_pe_2_nw[4][7]),
    .merge_valid_i_4_7                             (merge_valid_pe_2_nw[4][7]),
    .merge_ready_o_4_7                             (merge_ready_nw_2_pe[4][7]),
    .gather_data_i_4_7                             (gather_data_pe_2_nw[4][7]),
    .gather_valid_i_4_7                            (gather_valid_pe_2_nw[4][7]),
    .gather_ready_o_4_7                            (gather_ready_nw_2_pe[4][7]),

    .cast_data_o_4_7                               (cast_data_nw_2_pe[4][7]),
    .cast_valid_o_4_7                              (cast_valid_nw_2_pe[4][7]),
    .cast_ready_i_4_7                              (cast_ready_pe_2_nw[4][7]),
    .merge_data_o_4_7                              (merge_data_nw_2_pe[4][7]),
    .merge_valid_o_4_7                             (merge_valid_nw_2_pe[4][7]),
    .merge_ready_i_4_7                             (merge_ready_pe_2_nw[4][7]),
    .gather_data_o_4_7                             (gather_data_nw_2_pe[4][7]),
    .gather_valid_o_4_7                            (gather_valid_nw_2_pe[4][7]),
    .gather_ready_i_4_7                            (gather_ready_pe_2_nw[4][7]),
    .cast_data_i_4_8                               (cast_data_pe_2_nw[4][8]),
    .cast_valid_i_4_8                              (cast_valid_pe_2_nw[4][8]),
    .cast_ready_o_4_8                              (cast_ready_nw_2_pe[4][8]),
    .merge_data_i_4_8                              (merge_data_pe_2_nw[4][8]),
    .merge_valid_i_4_8                             (merge_valid_pe_2_nw[4][8]),
    .merge_ready_o_4_8                             (merge_ready_nw_2_pe[4][8]),
    .gather_data_i_4_8                             (gather_data_pe_2_nw[4][8]),
    .gather_valid_i_4_8                            (gather_valid_pe_2_nw[4][8]),
    .gather_ready_o_4_8                            (gather_ready_nw_2_pe[4][8]),

    .cast_data_o_4_8                               (cast_data_nw_2_pe[4][8]),
    .cast_valid_o_4_8                              (cast_valid_nw_2_pe[4][8]),
    .cast_ready_i_4_8                              (cast_ready_pe_2_nw[4][8]),
    .merge_data_o_4_8                              (merge_data_nw_2_pe[4][8]),
    .merge_valid_o_4_8                             (merge_valid_nw_2_pe[4][8]),
    .merge_ready_i_4_8                             (merge_ready_pe_2_nw[4][8]),
    .gather_data_o_4_8                             (gather_data_nw_2_pe[4][8]),
    .gather_valid_o_4_8                            (gather_valid_nw_2_pe[4][8]),
    .gather_ready_i_4_8                            (gather_ready_pe_2_nw[4][8]),
    .cast_data_i_4_9                               (cast_data_pe_2_nw[4][9]),
    .cast_valid_i_4_9                              (cast_valid_pe_2_nw[4][9]),
    .cast_ready_o_4_9                              (cast_ready_nw_2_pe[4][9]),
    .merge_data_i_4_9                              (merge_data_pe_2_nw[4][9]),
    .merge_valid_i_4_9                             (merge_valid_pe_2_nw[4][9]),
    .merge_ready_o_4_9                             (merge_ready_nw_2_pe[4][9]),
    .gather_data_i_4_9                             (gather_data_pe_2_nw[4][9]),
    .gather_valid_i_4_9                            (gather_valid_pe_2_nw[4][9]),
    .gather_ready_o_4_9                            (gather_ready_nw_2_pe[4][9]),

    .cast_data_o_4_9                               (cast_data_nw_2_pe[4][9]),
    .cast_valid_o_4_9                              (cast_valid_nw_2_pe[4][9]),
    .cast_ready_i_4_9                              (cast_ready_pe_2_nw[4][9]),
    .merge_data_o_4_9                              (merge_data_nw_2_pe[4][9]),
    .merge_valid_o_4_9                             (merge_valid_nw_2_pe[4][9]),
    .merge_ready_i_4_9                             (merge_ready_pe_2_nw[4][9]),
    .gather_data_o_4_9                             (gather_data_nw_2_pe[4][9]),
    .gather_valid_o_4_9                            (gather_valid_nw_2_pe[4][9]),
    .gather_ready_i_4_9                            (gather_ready_pe_2_nw[4][9])
);

virtual_pe #(
    .cast_out                                          (cast_out_0_0),
    .merge_in                                          (merge_in_0_0),
    .merge_out                                         (merge_out_0_0),
    .gather_in                                         (gather_in_0_0),
    .gather_out                                        (gather_out_0_0),
    .x                                                 (0),
    .y                                                 (0)
)vpe_0_0(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[0][0]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[0][0]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[0][0]),
    .cast_data_o                                       (cast_data_pe_2_nw[0][0]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[0][0]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[0][0]),
    .merge_data_i                                      (merge_data_nw_2_pe[0][0]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[0][0]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[0][0]),
    .merge_data_o                                      (merge_data_pe_2_nw[0][0]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[0][0]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[0][0]),
    .gather_data_i                                     (gather_data_nw_2_pe[0][0]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[0][0]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[0][0]),
    .gather_data_o                                     (gather_data_pe_2_nw[0][0]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[0][0]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[0][0])
);


virtual_pe #(
    .cast_out                                          (cast_out_0_1),
    .merge_in                                          (merge_in_0_1),
    .merge_out                                         (merge_out_0_1),
    .gather_in                                         (gather_in_0_1),
    .gather_out                                        (gather_out_0_1),
    .x                                                 (0),
    .y                                                 (1)
)vpe_0_1(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[0][1]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[0][1]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[0][1]),
    .cast_data_o                                       (cast_data_pe_2_nw[0][1]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[0][1]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[0][1]),
    .merge_data_i                                      (merge_data_nw_2_pe[0][1]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[0][1]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[0][1]),
    .merge_data_o                                      (merge_data_pe_2_nw[0][1]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[0][1]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[0][1]),
    .gather_data_i                                     (gather_data_nw_2_pe[0][1]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[0][1]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[0][1]),
    .gather_data_o                                     (gather_data_pe_2_nw[0][1]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[0][1]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[0][1])
);


virtual_pe #(
    .cast_out                                          (cast_out_0_2),
    .merge_in                                          (merge_in_0_2),
    .merge_out                                         (merge_out_0_2),
    .gather_in                                         (gather_in_0_2),
    .gather_out                                        (gather_out_0_2),
    .x                                                 (0),
    .y                                                 (2)
)vpe_0_2(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[0][2]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[0][2]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[0][2]),
    .cast_data_o                                       (cast_data_pe_2_nw[0][2]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[0][2]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[0][2]),
    .merge_data_i                                      (merge_data_nw_2_pe[0][2]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[0][2]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[0][2]),
    .merge_data_o                                      (merge_data_pe_2_nw[0][2]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[0][2]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[0][2]),
    .gather_data_i                                     (gather_data_nw_2_pe[0][2]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[0][2]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[0][2]),
    .gather_data_o                                     (gather_data_pe_2_nw[0][2]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[0][2]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[0][2])
);


virtual_pe #(
    .cast_out                                          (cast_out_0_3),
    .merge_in                                          (merge_in_0_3),
    .merge_out                                         (merge_out_0_3),
    .gather_in                                         (gather_in_0_3),
    .gather_out                                        (gather_out_0_3),
    .x                                                 (0),
    .y                                                 (3)
)vpe_0_3(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[0][3]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[0][3]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[0][3]),
    .cast_data_o                                       (cast_data_pe_2_nw[0][3]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[0][3]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[0][3]),
    .merge_data_i                                      (merge_data_nw_2_pe[0][3]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[0][3]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[0][3]),
    .merge_data_o                                      (merge_data_pe_2_nw[0][3]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[0][3]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[0][3]),
    .gather_data_i                                     (gather_data_nw_2_pe[0][3]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[0][3]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[0][3]),
    .gather_data_o                                     (gather_data_pe_2_nw[0][3]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[0][3]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[0][3])
);


virtual_pe #(
    .cast_out                                          (cast_out_0_4),
    .merge_in                                          (merge_in_0_4),
    .merge_out                                         (merge_out_0_4),
    .gather_in                                         (gather_in_0_4),
    .gather_out                                        (gather_out_0_4),
    .x                                                 (0),
    .y                                                 (4)
)vpe_0_4(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[0][4]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[0][4]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[0][4]),
    .cast_data_o                                       (cast_data_pe_2_nw[0][4]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[0][4]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[0][4]),
    .merge_data_i                                      (merge_data_nw_2_pe[0][4]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[0][4]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[0][4]),
    .merge_data_o                                      (merge_data_pe_2_nw[0][4]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[0][4]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[0][4]),
    .gather_data_i                                     (gather_data_nw_2_pe[0][4]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[0][4]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[0][4]),
    .gather_data_o                                     (gather_data_pe_2_nw[0][4]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[0][4]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[0][4])
);


virtual_pe #(
    .cast_out                                          (cast_out_0_5),
    .merge_in                                          (merge_in_0_5),
    .merge_out                                         (merge_out_0_5),
    .gather_in                                         (gather_in_0_5),
    .gather_out                                        (gather_out_0_5),
    .x                                                 (0),
    .y                                                 (5)
)vpe_0_5(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[0][5]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[0][5]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[0][5]),
    .cast_data_o                                       (cast_data_pe_2_nw[0][5]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[0][5]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[0][5]),
    .merge_data_i                                      (merge_data_nw_2_pe[0][5]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[0][5]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[0][5]),
    .merge_data_o                                      (merge_data_pe_2_nw[0][5]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[0][5]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[0][5]),
    .gather_data_i                                     (gather_data_nw_2_pe[0][5]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[0][5]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[0][5]),
    .gather_data_o                                     (gather_data_pe_2_nw[0][5]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[0][5]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[0][5])
);


virtual_pe #(
    .cast_out                                          (cast_out_0_6),
    .merge_in                                          (merge_in_0_6),
    .merge_out                                         (merge_out_0_6),
    .gather_in                                         (gather_in_0_6),
    .gather_out                                        (gather_out_0_6),
    .x                                                 (0),
    .y                                                 (6)
)vpe_0_6(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[0][6]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[0][6]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[0][6]),
    .cast_data_o                                       (cast_data_pe_2_nw[0][6]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[0][6]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[0][6]),
    .merge_data_i                                      (merge_data_nw_2_pe[0][6]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[0][6]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[0][6]),
    .merge_data_o                                      (merge_data_pe_2_nw[0][6]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[0][6]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[0][6]),
    .gather_data_i                                     (gather_data_nw_2_pe[0][6]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[0][6]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[0][6]),
    .gather_data_o                                     (gather_data_pe_2_nw[0][6]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[0][6]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[0][6])
);


virtual_pe #(
    .cast_out                                          (cast_out_0_7),
    .merge_in                                          (merge_in_0_7),
    .merge_out                                         (merge_out_0_7),
    .gather_in                                         (gather_in_0_7),
    .gather_out                                        (gather_out_0_7),
    .x                                                 (0),
    .y                                                 (7)
)vpe_0_7(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[0][7]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[0][7]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[0][7]),
    .cast_data_o                                       (cast_data_pe_2_nw[0][7]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[0][7]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[0][7]),
    .merge_data_i                                      (merge_data_nw_2_pe[0][7]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[0][7]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[0][7]),
    .merge_data_o                                      (merge_data_pe_2_nw[0][7]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[0][7]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[0][7]),
    .gather_data_i                                     (gather_data_nw_2_pe[0][7]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[0][7]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[0][7]),
    .gather_data_o                                     (gather_data_pe_2_nw[0][7]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[0][7]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[0][7])
);


virtual_pe #(
    .cast_out                                          (cast_out_0_8),
    .merge_in                                          (merge_in_0_8),
    .merge_out                                         (merge_out_0_8),
    .gather_in                                         (gather_in_0_8),
    .gather_out                                        (gather_out_0_8),
    .x                                                 (0),
    .y                                                 (8)
)vpe_0_8(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[0][8]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[0][8]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[0][8]),
    .cast_data_o                                       (cast_data_pe_2_nw[0][8]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[0][8]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[0][8]),
    .merge_data_i                                      (merge_data_nw_2_pe[0][8]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[0][8]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[0][8]),
    .merge_data_o                                      (merge_data_pe_2_nw[0][8]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[0][8]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[0][8]),
    .gather_data_i                                     (gather_data_nw_2_pe[0][8]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[0][8]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[0][8]),
    .gather_data_o                                     (gather_data_pe_2_nw[0][8]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[0][8]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[0][8])
);


virtual_pe #(
    .cast_out                                          (cast_out_0_9),
    .merge_in                                          (merge_in_0_9),
    .merge_out                                         (merge_out_0_9),
    .gather_in                                         (gather_in_0_9),
    .gather_out                                        (gather_out_0_9),
    .x                                                 (0),
    .y                                                 (9)
)vpe_0_9(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[0][9]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[0][9]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[0][9]),
    .cast_data_o                                       (cast_data_pe_2_nw[0][9]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[0][9]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[0][9]),
    .merge_data_i                                      (merge_data_nw_2_pe[0][9]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[0][9]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[0][9]),
    .merge_data_o                                      (merge_data_pe_2_nw[0][9]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[0][9]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[0][9]),
    .gather_data_i                                     (gather_data_nw_2_pe[0][9]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[0][9]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[0][9]),
    .gather_data_o                                     (gather_data_pe_2_nw[0][9]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[0][9]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[0][9])
);


virtual_pe #(
    .cast_out                                          (cast_out_1_0),
    .merge_in                                          (merge_in_1_0),
    .merge_out                                         (merge_out_1_0),
    .gather_in                                         (gather_in_1_0),
    .gather_out                                        (gather_out_1_0),
    .x                                                 (1),
    .y                                                 (0)
)vpe_1_0(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[1][0]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[1][0]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[1][0]),
    .cast_data_o                                       (cast_data_pe_2_nw[1][0]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[1][0]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[1][0]),
    .merge_data_i                                      (merge_data_nw_2_pe[1][0]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[1][0]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[1][0]),
    .merge_data_o                                      (merge_data_pe_2_nw[1][0]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[1][0]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[1][0]),
    .gather_data_i                                     (gather_data_nw_2_pe[1][0]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[1][0]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[1][0]),
    .gather_data_o                                     (gather_data_pe_2_nw[1][0]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[1][0]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[1][0])
);


virtual_pe #(
    .cast_out                                          (cast_out_1_1),
    .merge_in                                          (merge_in_1_1),
    .merge_out                                         (merge_out_1_1),
    .gather_in                                         (gather_in_1_1),
    .gather_out                                        (gather_out_1_1),
    .x                                                 (1),
    .y                                                 (1)
)vpe_1_1(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[1][1]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[1][1]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[1][1]),
    .cast_data_o                                       (cast_data_pe_2_nw[1][1]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[1][1]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[1][1]),
    .merge_data_i                                      (merge_data_nw_2_pe[1][1]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[1][1]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[1][1]),
    .merge_data_o                                      (merge_data_pe_2_nw[1][1]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[1][1]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[1][1]),
    .gather_data_i                                     (gather_data_nw_2_pe[1][1]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[1][1]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[1][1]),
    .gather_data_o                                     (gather_data_pe_2_nw[1][1]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[1][1]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[1][1])
);


virtual_pe #(
    .cast_out                                          (cast_out_1_2),
    .merge_in                                          (merge_in_1_2),
    .merge_out                                         (merge_out_1_2),
    .gather_in                                         (gather_in_1_2),
    .gather_out                                        (gather_out_1_2),
    .x                                                 (1),
    .y                                                 (2)
)vpe_1_2(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[1][2]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[1][2]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[1][2]),
    .cast_data_o                                       (cast_data_pe_2_nw[1][2]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[1][2]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[1][2]),
    .merge_data_i                                      (merge_data_nw_2_pe[1][2]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[1][2]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[1][2]),
    .merge_data_o                                      (merge_data_pe_2_nw[1][2]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[1][2]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[1][2]),
    .gather_data_i                                     (gather_data_nw_2_pe[1][2]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[1][2]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[1][2]),
    .gather_data_o                                     (gather_data_pe_2_nw[1][2]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[1][2]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[1][2])
);


virtual_pe #(
    .cast_out                                          (cast_out_1_3),
    .merge_in                                          (merge_in_1_3),
    .merge_out                                         (merge_out_1_3),
    .gather_in                                         (gather_in_1_3),
    .gather_out                                        (gather_out_1_3),
    .x                                                 (1),
    .y                                                 (3)
)vpe_1_3(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[1][3]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[1][3]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[1][3]),
    .cast_data_o                                       (cast_data_pe_2_nw[1][3]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[1][3]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[1][3]),
    .merge_data_i                                      (merge_data_nw_2_pe[1][3]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[1][3]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[1][3]),
    .merge_data_o                                      (merge_data_pe_2_nw[1][3]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[1][3]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[1][3]),
    .gather_data_i                                     (gather_data_nw_2_pe[1][3]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[1][3]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[1][3]),
    .gather_data_o                                     (gather_data_pe_2_nw[1][3]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[1][3]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[1][3])
);


virtual_pe #(
    .cast_out                                          (cast_out_1_4),
    .merge_in                                          (merge_in_1_4),
    .merge_out                                         (merge_out_1_4),
    .gather_in                                         (gather_in_1_4),
    .gather_out                                        (gather_out_1_4),
    .x                                                 (1),
    .y                                                 (4)
)vpe_1_4(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[1][4]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[1][4]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[1][4]),
    .cast_data_o                                       (cast_data_pe_2_nw[1][4]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[1][4]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[1][4]),
    .merge_data_i                                      (merge_data_nw_2_pe[1][4]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[1][4]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[1][4]),
    .merge_data_o                                      (merge_data_pe_2_nw[1][4]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[1][4]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[1][4]),
    .gather_data_i                                     (gather_data_nw_2_pe[1][4]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[1][4]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[1][4]),
    .gather_data_o                                     (gather_data_pe_2_nw[1][4]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[1][4]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[1][4])
);


virtual_pe #(
    .cast_out                                          (cast_out_1_5),
    .merge_in                                          (merge_in_1_5),
    .merge_out                                         (merge_out_1_5),
    .gather_in                                         (gather_in_1_5),
    .gather_out                                        (gather_out_1_5),
    .x                                                 (1),
    .y                                                 (5)
)vpe_1_5(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[1][5]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[1][5]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[1][5]),
    .cast_data_o                                       (cast_data_pe_2_nw[1][5]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[1][5]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[1][5]),
    .merge_data_i                                      (merge_data_nw_2_pe[1][5]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[1][5]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[1][5]),
    .merge_data_o                                      (merge_data_pe_2_nw[1][5]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[1][5]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[1][5]),
    .gather_data_i                                     (gather_data_nw_2_pe[1][5]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[1][5]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[1][5]),
    .gather_data_o                                     (gather_data_pe_2_nw[1][5]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[1][5]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[1][5])
);


virtual_pe #(
    .cast_out                                          (cast_out_1_6),
    .merge_in                                          (merge_in_1_6),
    .merge_out                                         (merge_out_1_6),
    .gather_in                                         (gather_in_1_6),
    .gather_out                                        (gather_out_1_6),
    .x                                                 (1),
    .y                                                 (6)
)vpe_1_6(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[1][6]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[1][6]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[1][6]),
    .cast_data_o                                       (cast_data_pe_2_nw[1][6]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[1][6]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[1][6]),
    .merge_data_i                                      (merge_data_nw_2_pe[1][6]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[1][6]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[1][6]),
    .merge_data_o                                      (merge_data_pe_2_nw[1][6]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[1][6]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[1][6]),
    .gather_data_i                                     (gather_data_nw_2_pe[1][6]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[1][6]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[1][6]),
    .gather_data_o                                     (gather_data_pe_2_nw[1][6]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[1][6]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[1][6])
);


virtual_pe #(
    .cast_out                                          (cast_out_1_7),
    .merge_in                                          (merge_in_1_7),
    .merge_out                                         (merge_out_1_7),
    .gather_in                                         (gather_in_1_7),
    .gather_out                                        (gather_out_1_7),
    .x                                                 (1),
    .y                                                 (7)
)vpe_1_7(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[1][7]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[1][7]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[1][7]),
    .cast_data_o                                       (cast_data_pe_2_nw[1][7]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[1][7]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[1][7]),
    .merge_data_i                                      (merge_data_nw_2_pe[1][7]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[1][7]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[1][7]),
    .merge_data_o                                      (merge_data_pe_2_nw[1][7]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[1][7]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[1][7]),
    .gather_data_i                                     (gather_data_nw_2_pe[1][7]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[1][7]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[1][7]),
    .gather_data_o                                     (gather_data_pe_2_nw[1][7]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[1][7]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[1][7])
);


virtual_pe #(
    .cast_out                                          (cast_out_1_8),
    .merge_in                                          (merge_in_1_8),
    .merge_out                                         (merge_out_1_8),
    .gather_in                                         (gather_in_1_8),
    .gather_out                                        (gather_out_1_8),
    .x                                                 (1),
    .y                                                 (8)
)vpe_1_8(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[1][8]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[1][8]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[1][8]),
    .cast_data_o                                       (cast_data_pe_2_nw[1][8]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[1][8]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[1][8]),
    .merge_data_i                                      (merge_data_nw_2_pe[1][8]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[1][8]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[1][8]),
    .merge_data_o                                      (merge_data_pe_2_nw[1][8]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[1][8]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[1][8]),
    .gather_data_i                                     (gather_data_nw_2_pe[1][8]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[1][8]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[1][8]),
    .gather_data_o                                     (gather_data_pe_2_nw[1][8]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[1][8]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[1][8])
);


virtual_pe #(
    .cast_out                                          (cast_out_1_9),
    .merge_in                                          (merge_in_1_9),
    .merge_out                                         (merge_out_1_9),
    .gather_in                                         (gather_in_1_9),
    .gather_out                                        (gather_out_1_9),
    .x                                                 (1),
    .y                                                 (9)
)vpe_1_9(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[1][9]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[1][9]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[1][9]),
    .cast_data_o                                       (cast_data_pe_2_nw[1][9]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[1][9]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[1][9]),
    .merge_data_i                                      (merge_data_nw_2_pe[1][9]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[1][9]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[1][9]),
    .merge_data_o                                      (merge_data_pe_2_nw[1][9]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[1][9]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[1][9]),
    .gather_data_i                                     (gather_data_nw_2_pe[1][9]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[1][9]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[1][9]),
    .gather_data_o                                     (gather_data_pe_2_nw[1][9]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[1][9]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[1][9])
);


virtual_pe #(
    .cast_out                                          (cast_out_2_0),
    .merge_in                                          (merge_in_2_0),
    .merge_out                                         (merge_out_2_0),
    .gather_in                                         (gather_in_2_0),
    .gather_out                                        (gather_out_2_0),
    .x                                                 (2),
    .y                                                 (0)
)vpe_2_0(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[2][0]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[2][0]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[2][0]),
    .cast_data_o                                       (cast_data_pe_2_nw[2][0]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[2][0]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[2][0]),
    .merge_data_i                                      (merge_data_nw_2_pe[2][0]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[2][0]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[2][0]),
    .merge_data_o                                      (merge_data_pe_2_nw[2][0]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[2][0]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[2][0]),
    .gather_data_i                                     (gather_data_nw_2_pe[2][0]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[2][0]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[2][0]),
    .gather_data_o                                     (gather_data_pe_2_nw[2][0]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[2][0]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[2][0])
);


virtual_pe #(
    .cast_out                                          (cast_out_2_1),
    .merge_in                                          (merge_in_2_1),
    .merge_out                                         (merge_out_2_1),
    .gather_in                                         (gather_in_2_1),
    .gather_out                                        (gather_out_2_1),
    .x                                                 (2),
    .y                                                 (1)
)vpe_2_1(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[2][1]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[2][1]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[2][1]),
    .cast_data_o                                       (cast_data_pe_2_nw[2][1]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[2][1]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[2][1]),
    .merge_data_i                                      (merge_data_nw_2_pe[2][1]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[2][1]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[2][1]),
    .merge_data_o                                      (merge_data_pe_2_nw[2][1]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[2][1]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[2][1]),
    .gather_data_i                                     (gather_data_nw_2_pe[2][1]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[2][1]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[2][1]),
    .gather_data_o                                     (gather_data_pe_2_nw[2][1]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[2][1]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[2][1])
);


virtual_pe #(
    .cast_out                                          (cast_out_2_2),
    .merge_in                                          (merge_in_2_2),
    .merge_out                                         (merge_out_2_2),
    .gather_in                                         (gather_in_2_2),
    .gather_out                                        (gather_out_2_2),
    .x                                                 (2),
    .y                                                 (2)
)vpe_2_2(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[2][2]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[2][2]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[2][2]),
    .cast_data_o                                       (cast_data_pe_2_nw[2][2]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[2][2]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[2][2]),
    .merge_data_i                                      (merge_data_nw_2_pe[2][2]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[2][2]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[2][2]),
    .merge_data_o                                      (merge_data_pe_2_nw[2][2]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[2][2]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[2][2]),
    .gather_data_i                                     (gather_data_nw_2_pe[2][2]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[2][2]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[2][2]),
    .gather_data_o                                     (gather_data_pe_2_nw[2][2]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[2][2]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[2][2])
);


virtual_pe #(
    .cast_out                                          (cast_out_2_3),
    .merge_in                                          (merge_in_2_3),
    .merge_out                                         (merge_out_2_3),
    .gather_in                                         (gather_in_2_3),
    .gather_out                                        (gather_out_2_3),
    .x                                                 (2),
    .y                                                 (3)
)vpe_2_3(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[2][3]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[2][3]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[2][3]),
    .cast_data_o                                       (cast_data_pe_2_nw[2][3]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[2][3]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[2][3]),
    .merge_data_i                                      (merge_data_nw_2_pe[2][3]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[2][3]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[2][3]),
    .merge_data_o                                      (merge_data_pe_2_nw[2][3]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[2][3]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[2][3]),
    .gather_data_i                                     (gather_data_nw_2_pe[2][3]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[2][3]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[2][3]),
    .gather_data_o                                     (gather_data_pe_2_nw[2][3]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[2][3]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[2][3])
);


virtual_pe #(
    .cast_out                                          (cast_out_2_4),
    .merge_in                                          (merge_in_2_4),
    .merge_out                                         (merge_out_2_4),
    .gather_in                                         (gather_in_2_4),
    .gather_out                                        (gather_out_2_4),
    .x                                                 (2),
    .y                                                 (4)
)vpe_2_4(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[2][4]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[2][4]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[2][4]),
    .cast_data_o                                       (cast_data_pe_2_nw[2][4]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[2][4]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[2][4]),
    .merge_data_i                                      (merge_data_nw_2_pe[2][4]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[2][4]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[2][4]),
    .merge_data_o                                      (merge_data_pe_2_nw[2][4]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[2][4]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[2][4]),
    .gather_data_i                                     (gather_data_nw_2_pe[2][4]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[2][4]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[2][4]),
    .gather_data_o                                     (gather_data_pe_2_nw[2][4]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[2][4]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[2][4])
);


virtual_pe #(
    .cast_out                                          (cast_out_2_5),
    .merge_in                                          (merge_in_2_5),
    .merge_out                                         (merge_out_2_5),
    .gather_in                                         (gather_in_2_5),
    .gather_out                                        (gather_out_2_5),
    .x                                                 (2),
    .y                                                 (5)
)vpe_2_5(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[2][5]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[2][5]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[2][5]),
    .cast_data_o                                       (cast_data_pe_2_nw[2][5]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[2][5]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[2][5]),
    .merge_data_i                                      (merge_data_nw_2_pe[2][5]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[2][5]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[2][5]),
    .merge_data_o                                      (merge_data_pe_2_nw[2][5]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[2][5]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[2][5]),
    .gather_data_i                                     (gather_data_nw_2_pe[2][5]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[2][5]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[2][5]),
    .gather_data_o                                     (gather_data_pe_2_nw[2][5]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[2][5]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[2][5])
);


virtual_pe #(
    .cast_out                                          (cast_out_2_6),
    .merge_in                                          (merge_in_2_6),
    .merge_out                                         (merge_out_2_6),
    .gather_in                                         (gather_in_2_6),
    .gather_out                                        (gather_out_2_6),
    .x                                                 (2),
    .y                                                 (6)
)vpe_2_6(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[2][6]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[2][6]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[2][6]),
    .cast_data_o                                       (cast_data_pe_2_nw[2][6]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[2][6]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[2][6]),
    .merge_data_i                                      (merge_data_nw_2_pe[2][6]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[2][6]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[2][6]),
    .merge_data_o                                      (merge_data_pe_2_nw[2][6]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[2][6]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[2][6]),
    .gather_data_i                                     (gather_data_nw_2_pe[2][6]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[2][6]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[2][6]),
    .gather_data_o                                     (gather_data_pe_2_nw[2][6]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[2][6]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[2][6])
);


virtual_pe #(
    .cast_out                                          (cast_out_2_7),
    .merge_in                                          (merge_in_2_7),
    .merge_out                                         (merge_out_2_7),
    .gather_in                                         (gather_in_2_7),
    .gather_out                                        (gather_out_2_7),
    .x                                                 (2),
    .y                                                 (7)
)vpe_2_7(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[2][7]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[2][7]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[2][7]),
    .cast_data_o                                       (cast_data_pe_2_nw[2][7]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[2][7]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[2][7]),
    .merge_data_i                                      (merge_data_nw_2_pe[2][7]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[2][7]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[2][7]),
    .merge_data_o                                      (merge_data_pe_2_nw[2][7]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[2][7]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[2][7]),
    .gather_data_i                                     (gather_data_nw_2_pe[2][7]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[2][7]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[2][7]),
    .gather_data_o                                     (gather_data_pe_2_nw[2][7]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[2][7]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[2][7])
);


virtual_pe #(
    .cast_out                                          (cast_out_2_8),
    .merge_in                                          (merge_in_2_8),
    .merge_out                                         (merge_out_2_8),
    .gather_in                                         (gather_in_2_8),
    .gather_out                                        (gather_out_2_8),
    .x                                                 (2),
    .y                                                 (8)
)vpe_2_8(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[2][8]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[2][8]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[2][8]),
    .cast_data_o                                       (cast_data_pe_2_nw[2][8]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[2][8]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[2][8]),
    .merge_data_i                                      (merge_data_nw_2_pe[2][8]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[2][8]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[2][8]),
    .merge_data_o                                      (merge_data_pe_2_nw[2][8]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[2][8]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[2][8]),
    .gather_data_i                                     (gather_data_nw_2_pe[2][8]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[2][8]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[2][8]),
    .gather_data_o                                     (gather_data_pe_2_nw[2][8]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[2][8]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[2][8])
);


virtual_pe #(
    .cast_out                                          (cast_out_2_9),
    .merge_in                                          (merge_in_2_9),
    .merge_out                                         (merge_out_2_9),
    .gather_in                                         (gather_in_2_9),
    .gather_out                                        (gather_out_2_9),
    .x                                                 (2),
    .y                                                 (9)
)vpe_2_9(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[2][9]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[2][9]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[2][9]),
    .cast_data_o                                       (cast_data_pe_2_nw[2][9]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[2][9]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[2][9]),
    .merge_data_i                                      (merge_data_nw_2_pe[2][9]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[2][9]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[2][9]),
    .merge_data_o                                      (merge_data_pe_2_nw[2][9]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[2][9]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[2][9]),
    .gather_data_i                                     (gather_data_nw_2_pe[2][9]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[2][9]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[2][9]),
    .gather_data_o                                     (gather_data_pe_2_nw[2][9]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[2][9]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[2][9])
);


virtual_pe #(
    .cast_out                                          (cast_out_3_0),
    .merge_in                                          (merge_in_3_0),
    .merge_out                                         (merge_out_3_0),
    .gather_in                                         (gather_in_3_0),
    .gather_out                                        (gather_out_3_0),
    .x                                                 (3),
    .y                                                 (0)
)vpe_3_0(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[3][0]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[3][0]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[3][0]),
    .cast_data_o                                       (cast_data_pe_2_nw[3][0]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[3][0]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[3][0]),
    .merge_data_i                                      (merge_data_nw_2_pe[3][0]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[3][0]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[3][0]),
    .merge_data_o                                      (merge_data_pe_2_nw[3][0]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[3][0]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[3][0]),
    .gather_data_i                                     (gather_data_nw_2_pe[3][0]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[3][0]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[3][0]),
    .gather_data_o                                     (gather_data_pe_2_nw[3][0]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[3][0]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[3][0])
);


virtual_pe #(
    .cast_out                                          (cast_out_3_1),
    .merge_in                                          (merge_in_3_1),
    .merge_out                                         (merge_out_3_1),
    .gather_in                                         (gather_in_3_1),
    .gather_out                                        (gather_out_3_1),
    .x                                                 (3),
    .y                                                 (1)
)vpe_3_1(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[3][1]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[3][1]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[3][1]),
    .cast_data_o                                       (cast_data_pe_2_nw[3][1]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[3][1]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[3][1]),
    .merge_data_i                                      (merge_data_nw_2_pe[3][1]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[3][1]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[3][1]),
    .merge_data_o                                      (merge_data_pe_2_nw[3][1]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[3][1]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[3][1]),
    .gather_data_i                                     (gather_data_nw_2_pe[3][1]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[3][1]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[3][1]),
    .gather_data_o                                     (gather_data_pe_2_nw[3][1]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[3][1]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[3][1])
);


virtual_pe #(
    .cast_out                                          (cast_out_3_2),
    .merge_in                                          (merge_in_3_2),
    .merge_out                                         (merge_out_3_2),
    .gather_in                                         (gather_in_3_2),
    .gather_out                                        (gather_out_3_2),
    .x                                                 (3),
    .y                                                 (2)
)vpe_3_2(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[3][2]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[3][2]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[3][2]),
    .cast_data_o                                       (cast_data_pe_2_nw[3][2]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[3][2]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[3][2]),
    .merge_data_i                                      (merge_data_nw_2_pe[3][2]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[3][2]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[3][2]),
    .merge_data_o                                      (merge_data_pe_2_nw[3][2]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[3][2]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[3][2]),
    .gather_data_i                                     (gather_data_nw_2_pe[3][2]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[3][2]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[3][2]),
    .gather_data_o                                     (gather_data_pe_2_nw[3][2]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[3][2]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[3][2])
);


virtual_pe #(
    .cast_out                                          (cast_out_3_3),
    .merge_in                                          (merge_in_3_3),
    .merge_out                                         (merge_out_3_3),
    .gather_in                                         (gather_in_3_3),
    .gather_out                                        (gather_out_3_3),
    .x                                                 (3),
    .y                                                 (3)
)vpe_3_3(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[3][3]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[3][3]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[3][3]),
    .cast_data_o                                       (cast_data_pe_2_nw[3][3]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[3][3]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[3][3]),
    .merge_data_i                                      (merge_data_nw_2_pe[3][3]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[3][3]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[3][3]),
    .merge_data_o                                      (merge_data_pe_2_nw[3][3]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[3][3]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[3][3]),
    .gather_data_i                                     (gather_data_nw_2_pe[3][3]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[3][3]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[3][3]),
    .gather_data_o                                     (gather_data_pe_2_nw[3][3]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[3][3]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[3][3])
);


virtual_pe #(
    .cast_out                                          (cast_out_3_4),
    .merge_in                                          (merge_in_3_4),
    .merge_out                                         (merge_out_3_4),
    .gather_in                                         (gather_in_3_4),
    .gather_out                                        (gather_out_3_4),
    .x                                                 (3),
    .y                                                 (4)
)vpe_3_4(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[3][4]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[3][4]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[3][4]),
    .cast_data_o                                       (cast_data_pe_2_nw[3][4]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[3][4]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[3][4]),
    .merge_data_i                                      (merge_data_nw_2_pe[3][4]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[3][4]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[3][4]),
    .merge_data_o                                      (merge_data_pe_2_nw[3][4]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[3][4]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[3][4]),
    .gather_data_i                                     (gather_data_nw_2_pe[3][4]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[3][4]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[3][4]),
    .gather_data_o                                     (gather_data_pe_2_nw[3][4]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[3][4]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[3][4])
);


virtual_pe #(
    .cast_out                                          (cast_out_3_5),
    .merge_in                                          (merge_in_3_5),
    .merge_out                                         (merge_out_3_5),
    .gather_in                                         (gather_in_3_5),
    .gather_out                                        (gather_out_3_5),
    .x                                                 (3),
    .y                                                 (5)
)vpe_3_5(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[3][5]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[3][5]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[3][5]),
    .cast_data_o                                       (cast_data_pe_2_nw[3][5]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[3][5]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[3][5]),
    .merge_data_i                                      (merge_data_nw_2_pe[3][5]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[3][5]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[3][5]),
    .merge_data_o                                      (merge_data_pe_2_nw[3][5]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[3][5]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[3][5]),
    .gather_data_i                                     (gather_data_nw_2_pe[3][5]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[3][5]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[3][5]),
    .gather_data_o                                     (gather_data_pe_2_nw[3][5]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[3][5]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[3][5])
);


virtual_pe #(
    .cast_out                                          (cast_out_3_6),
    .merge_in                                          (merge_in_3_6),
    .merge_out                                         (merge_out_3_6),
    .gather_in                                         (gather_in_3_6),
    .gather_out                                        (gather_out_3_6),
    .x                                                 (3),
    .y                                                 (6)
)vpe_3_6(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[3][6]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[3][6]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[3][6]),
    .cast_data_o                                       (cast_data_pe_2_nw[3][6]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[3][6]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[3][6]),
    .merge_data_i                                      (merge_data_nw_2_pe[3][6]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[3][6]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[3][6]),
    .merge_data_o                                      (merge_data_pe_2_nw[3][6]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[3][6]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[3][6]),
    .gather_data_i                                     (gather_data_nw_2_pe[3][6]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[3][6]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[3][6]),
    .gather_data_o                                     (gather_data_pe_2_nw[3][6]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[3][6]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[3][6])
);


virtual_pe #(
    .cast_out                                          (cast_out_3_7),
    .merge_in                                          (merge_in_3_7),
    .merge_out                                         (merge_out_3_7),
    .gather_in                                         (gather_in_3_7),
    .gather_out                                        (gather_out_3_7),
    .x                                                 (3),
    .y                                                 (7)
)vpe_3_7(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[3][7]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[3][7]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[3][7]),
    .cast_data_o                                       (cast_data_pe_2_nw[3][7]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[3][7]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[3][7]),
    .merge_data_i                                      (merge_data_nw_2_pe[3][7]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[3][7]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[3][7]),
    .merge_data_o                                      (merge_data_pe_2_nw[3][7]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[3][7]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[3][7]),
    .gather_data_i                                     (gather_data_nw_2_pe[3][7]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[3][7]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[3][7]),
    .gather_data_o                                     (gather_data_pe_2_nw[3][7]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[3][7]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[3][7])
);


virtual_pe #(
    .cast_out                                          (cast_out_3_8),
    .merge_in                                          (merge_in_3_8),
    .merge_out                                         (merge_out_3_8),
    .gather_in                                         (gather_in_3_8),
    .gather_out                                        (gather_out_3_8),
    .x                                                 (3),
    .y                                                 (8)
)vpe_3_8(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[3][8]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[3][8]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[3][8]),
    .cast_data_o                                       (cast_data_pe_2_nw[3][8]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[3][8]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[3][8]),
    .merge_data_i                                      (merge_data_nw_2_pe[3][8]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[3][8]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[3][8]),
    .merge_data_o                                      (merge_data_pe_2_nw[3][8]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[3][8]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[3][8]),
    .gather_data_i                                     (gather_data_nw_2_pe[3][8]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[3][8]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[3][8]),
    .gather_data_o                                     (gather_data_pe_2_nw[3][8]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[3][8]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[3][8])
);


virtual_pe #(
    .cast_out                                          (cast_out_3_9),
    .merge_in                                          (merge_in_3_9),
    .merge_out                                         (merge_out_3_9),
    .gather_in                                         (gather_in_3_9),
    .gather_out                                        (gather_out_3_9),
    .x                                                 (3),
    .y                                                 (9)
)vpe_3_9(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[3][9]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[3][9]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[3][9]),
    .cast_data_o                                       (cast_data_pe_2_nw[3][9]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[3][9]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[3][9]),
    .merge_data_i                                      (merge_data_nw_2_pe[3][9]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[3][9]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[3][9]),
    .merge_data_o                                      (merge_data_pe_2_nw[3][9]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[3][9]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[3][9]),
    .gather_data_i                                     (gather_data_nw_2_pe[3][9]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[3][9]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[3][9]),
    .gather_data_o                                     (gather_data_pe_2_nw[3][9]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[3][9]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[3][9])
);


virtual_pe #(
    .cast_out                                          (cast_out_4_0),
    .merge_in                                          (merge_in_4_0),
    .merge_out                                         (merge_out_4_0),
    .gather_in                                         (gather_in_4_0),
    .gather_out                                        (gather_out_4_0),
    .x                                                 (4),
    .y                                                 (0)
)vpe_4_0(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[4][0]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[4][0]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[4][0]),
    .cast_data_o                                       (cast_data_pe_2_nw[4][0]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[4][0]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[4][0]),
    .merge_data_i                                      (merge_data_nw_2_pe[4][0]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[4][0]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[4][0]),
    .merge_data_o                                      (merge_data_pe_2_nw[4][0]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[4][0]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[4][0]),
    .gather_data_i                                     (gather_data_nw_2_pe[4][0]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[4][0]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[4][0]),
    .gather_data_o                                     (gather_data_pe_2_nw[4][0]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[4][0]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[4][0])
);


virtual_pe #(
    .cast_out                                          (cast_out_4_1),
    .merge_in                                          (merge_in_4_1),
    .merge_out                                         (merge_out_4_1),
    .gather_in                                         (gather_in_4_1),
    .gather_out                                        (gather_out_4_1),
    .x                                                 (4),
    .y                                                 (1)
)vpe_4_1(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[4][1]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[4][1]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[4][1]),
    .cast_data_o                                       (cast_data_pe_2_nw[4][1]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[4][1]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[4][1]),
    .merge_data_i                                      (merge_data_nw_2_pe[4][1]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[4][1]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[4][1]),
    .merge_data_o                                      (merge_data_pe_2_nw[4][1]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[4][1]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[4][1]),
    .gather_data_i                                     (gather_data_nw_2_pe[4][1]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[4][1]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[4][1]),
    .gather_data_o                                     (gather_data_pe_2_nw[4][1]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[4][1]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[4][1])
);


virtual_pe #(
    .cast_out                                          (cast_out_4_2),
    .merge_in                                          (merge_in_4_2),
    .merge_out                                         (merge_out_4_2),
    .gather_in                                         (gather_in_4_2),
    .gather_out                                        (gather_out_4_2),
    .x                                                 (4),
    .y                                                 (2)
)vpe_4_2(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[4][2]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[4][2]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[4][2]),
    .cast_data_o                                       (cast_data_pe_2_nw[4][2]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[4][2]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[4][2]),
    .merge_data_i                                      (merge_data_nw_2_pe[4][2]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[4][2]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[4][2]),
    .merge_data_o                                      (merge_data_pe_2_nw[4][2]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[4][2]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[4][2]),
    .gather_data_i                                     (gather_data_nw_2_pe[4][2]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[4][2]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[4][2]),
    .gather_data_o                                     (gather_data_pe_2_nw[4][2]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[4][2]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[4][2])
);


virtual_pe #(
    .cast_out                                          (cast_out_4_3),
    .merge_in                                          (merge_in_4_3),
    .merge_out                                         (merge_out_4_3),
    .gather_in                                         (gather_in_4_3),
    .gather_out                                        (gather_out_4_3),
    .x                                                 (4),
    .y                                                 (3)
)vpe_4_3(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[4][3]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[4][3]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[4][3]),
    .cast_data_o                                       (cast_data_pe_2_nw[4][3]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[4][3]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[4][3]),
    .merge_data_i                                      (merge_data_nw_2_pe[4][3]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[4][3]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[4][3]),
    .merge_data_o                                      (merge_data_pe_2_nw[4][3]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[4][3]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[4][3]),
    .gather_data_i                                     (gather_data_nw_2_pe[4][3]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[4][3]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[4][3]),
    .gather_data_o                                     (gather_data_pe_2_nw[4][3]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[4][3]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[4][3])
);


virtual_pe #(
    .cast_out                                          (cast_out_4_4),
    .merge_in                                          (merge_in_4_4),
    .merge_out                                         (merge_out_4_4),
    .gather_in                                         (gather_in_4_4),
    .gather_out                                        (gather_out_4_4),
    .x                                                 (4),
    .y                                                 (4)
)vpe_4_4(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[4][4]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[4][4]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[4][4]),
    .cast_data_o                                       (cast_data_pe_2_nw[4][4]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[4][4]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[4][4]),
    .merge_data_i                                      (merge_data_nw_2_pe[4][4]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[4][4]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[4][4]),
    .merge_data_o                                      (merge_data_pe_2_nw[4][4]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[4][4]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[4][4]),
    .gather_data_i                                     (gather_data_nw_2_pe[4][4]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[4][4]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[4][4]),
    .gather_data_o                                     (gather_data_pe_2_nw[4][4]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[4][4]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[4][4])
);


virtual_pe #(
    .cast_out                                          (cast_out_4_5),
    .merge_in                                          (merge_in_4_5),
    .merge_out                                         (merge_out_4_5),
    .gather_in                                         (gather_in_4_5),
    .gather_out                                        (gather_out_4_5),
    .x                                                 (4),
    .y                                                 (5)
)vpe_4_5(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[4][5]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[4][5]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[4][5]),
    .cast_data_o                                       (cast_data_pe_2_nw[4][5]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[4][5]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[4][5]),
    .merge_data_i                                      (merge_data_nw_2_pe[4][5]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[4][5]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[4][5]),
    .merge_data_o                                      (merge_data_pe_2_nw[4][5]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[4][5]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[4][5]),
    .gather_data_i                                     (gather_data_nw_2_pe[4][5]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[4][5]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[4][5]),
    .gather_data_o                                     (gather_data_pe_2_nw[4][5]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[4][5]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[4][5])
);


virtual_pe #(
    .cast_out                                          (cast_out_4_6),
    .merge_in                                          (merge_in_4_6),
    .merge_out                                         (merge_out_4_6),
    .gather_in                                         (gather_in_4_6),
    .gather_out                                        (gather_out_4_6),
    .x                                                 (4),
    .y                                                 (6)
)vpe_4_6(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[4][6]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[4][6]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[4][6]),
    .cast_data_o                                       (cast_data_pe_2_nw[4][6]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[4][6]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[4][6]),
    .merge_data_i                                      (merge_data_nw_2_pe[4][6]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[4][6]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[4][6]),
    .merge_data_o                                      (merge_data_pe_2_nw[4][6]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[4][6]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[4][6]),
    .gather_data_i                                     (gather_data_nw_2_pe[4][6]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[4][6]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[4][6]),
    .gather_data_o                                     (gather_data_pe_2_nw[4][6]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[4][6]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[4][6])
);


virtual_pe #(
    .cast_out                                          (cast_out_4_7),
    .merge_in                                          (merge_in_4_7),
    .merge_out                                         (merge_out_4_7),
    .gather_in                                         (gather_in_4_7),
    .gather_out                                        (gather_out_4_7),
    .x                                                 (4),
    .y                                                 (7)
)vpe_4_7(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[4][7]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[4][7]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[4][7]),
    .cast_data_o                                       (cast_data_pe_2_nw[4][7]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[4][7]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[4][7]),
    .merge_data_i                                      (merge_data_nw_2_pe[4][7]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[4][7]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[4][7]),
    .merge_data_o                                      (merge_data_pe_2_nw[4][7]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[4][7]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[4][7]),
    .gather_data_i                                     (gather_data_nw_2_pe[4][7]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[4][7]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[4][7]),
    .gather_data_o                                     (gather_data_pe_2_nw[4][7]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[4][7]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[4][7])
);


virtual_pe #(
    .cast_out                                          (cast_out_4_8),
    .merge_in                                          (merge_in_4_8),
    .merge_out                                         (merge_out_4_8),
    .gather_in                                         (gather_in_4_8),
    .gather_out                                        (gather_out_4_8),
    .x                                                 (4),
    .y                                                 (8)
)vpe_4_8(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[4][8]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[4][8]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[4][8]),
    .cast_data_o                                       (cast_data_pe_2_nw[4][8]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[4][8]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[4][8]),
    .merge_data_i                                      (merge_data_nw_2_pe[4][8]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[4][8]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[4][8]),
    .merge_data_o                                      (merge_data_pe_2_nw[4][8]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[4][8]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[4][8]),
    .gather_data_i                                     (gather_data_nw_2_pe[4][8]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[4][8]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[4][8]),
    .gather_data_o                                     (gather_data_pe_2_nw[4][8]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[4][8]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[4][8])
);


virtual_pe #(
    .cast_out                                          (cast_out_4_9),
    .merge_in                                          (merge_in_4_9),
    .merge_out                                         (merge_out_4_9),
    .gather_in                                         (gather_in_4_9),
    .gather_out                                        (gather_out_4_9),
    .x                                                 (4),
    .y                                                 (9)
)vpe_4_9(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[4][9]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[4][9]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[4][9]),
    .cast_data_o                                       (cast_data_pe_2_nw[4][9]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[4][9]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[4][9]),
    .merge_data_i                                      (merge_data_nw_2_pe[4][9]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[4][9]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[4][9]),
    .merge_data_o                                      (merge_data_pe_2_nw[4][9]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[4][9]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[4][9]),
    .gather_data_i                                     (gather_data_nw_2_pe[4][9]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[4][9]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[4][9]),
    .gather_data_o                                     (gather_data_pe_2_nw[4][9]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[4][9]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[4][9])
);

endmodule
