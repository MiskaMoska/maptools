
//Cast Network
//Width: 10
//Height:25
`include "params.svh"
`include "cast_network_config.svh"

module cast_network(
    input       wire                            clk,
    input       wire                            rstn,

    //router local ports
    input       wire        [`DW-1:0]           data_i[`NOC_WIDTH][`NOC_HEIGHT],
    input       wire                            valid_i[`NOC_WIDTH][`NOC_HEIGHT],
    output      wire                            ready_o[`NOC_WIDTH][`NOC_HEIGHT],

    output      wire        [`DW-1:0]           data_o[`NOC_WIDTH][`NOC_HEIGHT],
    output      wire                            valid_o[`NOC_WIDTH][`NOC_HEIGHT],
    input       wire                            ready_i[`NOC_WIDTH][`NOC_HEIGHT],

    input       wire        [`DW-1:0]           data_i_stab,
    input       wire                            valid_i_stab,
    output      wire                            ready_o_stab,

    output      wire        [`DW-1:0]           data_o_flee0,
    output      wire                            valid_o_flee0,
    input       wire                            ready_i_flee0,

    output      wire        [`DW-1:0]           data_o_flee1,
    output      wire                            valid_o_flee1,
    input       wire                            ready_i_flee1,

    output      wire        [`DW-1:0]           data_o_flee2,
    output      wire                            valid_o_flee2,
    input       wire                            ready_i_flee2,

    output      wire        [`DW-1:0]           data_o_flee3,
    output      wire                            valid_o_flee3,
    input       wire                            ready_i_flee3,

    output      wire        [`DW-1:0]           data_o_flee4,
    output      wire                            valid_o_flee4,
    input       wire                            ready_i_flee4,

    output      wire        [`DW-1:0]           data_o_flee5,
    output      wire                            valid_o_flee5,
    input       wire                            ready_i_flee5,

    output      wire        [`DW-1:0]           data_o_flee6,
    output      wire                            valid_o_flee6,
    input       wire                            ready_i_flee6,

    output      wire        [`DW-1:0]           data_o_flee7,
    output      wire                            valid_o_flee7,
    input       wire                            ready_i_flee7,

    //credit update signal input
    input       wire                            credit_upd[`NOC_WIDTH][`NOC_HEIGHT]

);

//horizontal signals
wire    [`DW-1:0]   data_0_to_1,	data_1_to_0;
wire                valid_0_to_1,	valid_1_to_0;
wire                ready_0_to_1,	ready_1_to_0;
wire    [`DW-1:0]   data_1_to_2,	data_2_to_1;
wire                valid_1_to_2,	valid_2_to_1;
wire                ready_1_to_2,	ready_2_to_1;
wire    [`DW-1:0]   data_2_to_3,	data_3_to_2;
wire                valid_2_to_3,	valid_3_to_2;
wire                ready_2_to_3,	ready_3_to_2;
wire    [`DW-1:0]   data_3_to_4,	data_4_to_3;
wire                valid_3_to_4,	valid_4_to_3;
wire                ready_3_to_4,	ready_4_to_3;
wire    [`DW-1:0]   data_4_to_5,	data_5_to_4;
wire                valid_4_to_5,	valid_5_to_4;
wire                ready_4_to_5,	ready_5_to_4;
wire    [`DW-1:0]   data_5_to_6,	data_6_to_5;
wire                valid_5_to_6,	valid_6_to_5;
wire                ready_5_to_6,	ready_6_to_5;
wire    [`DW-1:0]   data_6_to_7,	data_7_to_6;
wire                valid_6_to_7,	valid_7_to_6;
wire                ready_6_to_7,	ready_7_to_6;
wire    [`DW-1:0]   data_7_to_8,	data_8_to_7;
wire                valid_7_to_8,	valid_8_to_7;
wire                ready_7_to_8,	ready_8_to_7;
wire    [`DW-1:0]   data_8_to_9,	data_9_to_8;
wire                valid_8_to_9,	valid_9_to_8;
wire                ready_8_to_9,	ready_9_to_8;
wire    [`DW-1:0]   data_10_to_11,	data_11_to_10;
wire                valid_10_to_11,	valid_11_to_10;
wire                ready_10_to_11,	ready_11_to_10;
wire    [`DW-1:0]   data_11_to_12,	data_12_to_11;
wire                valid_11_to_12,	valid_12_to_11;
wire                ready_11_to_12,	ready_12_to_11;
wire    [`DW-1:0]   data_12_to_13,	data_13_to_12;
wire                valid_12_to_13,	valid_13_to_12;
wire                ready_12_to_13,	ready_13_to_12;
wire    [`DW-1:0]   data_13_to_14,	data_14_to_13;
wire                valid_13_to_14,	valid_14_to_13;
wire                ready_13_to_14,	ready_14_to_13;
wire    [`DW-1:0]   data_14_to_15,	data_15_to_14;
wire                valid_14_to_15,	valid_15_to_14;
wire                ready_14_to_15,	ready_15_to_14;
wire    [`DW-1:0]   data_15_to_16,	data_16_to_15;
wire                valid_15_to_16,	valid_16_to_15;
wire                ready_15_to_16,	ready_16_to_15;
wire    [`DW-1:0]   data_16_to_17,	data_17_to_16;
wire                valid_16_to_17,	valid_17_to_16;
wire                ready_16_to_17,	ready_17_to_16;
wire    [`DW-1:0]   data_17_to_18,	data_18_to_17;
wire                valid_17_to_18,	valid_18_to_17;
wire                ready_17_to_18,	ready_18_to_17;
wire    [`DW-1:0]   data_18_to_19,	data_19_to_18;
wire                valid_18_to_19,	valid_19_to_18;
wire                ready_18_to_19,	ready_19_to_18;
wire    [`DW-1:0]   data_20_to_21,	data_21_to_20;
wire                valid_20_to_21,	valid_21_to_20;
wire                ready_20_to_21,	ready_21_to_20;
wire    [`DW-1:0]   data_21_to_22,	data_22_to_21;
wire                valid_21_to_22,	valid_22_to_21;
wire                ready_21_to_22,	ready_22_to_21;
wire    [`DW-1:0]   data_22_to_23,	data_23_to_22;
wire                valid_22_to_23,	valid_23_to_22;
wire                ready_22_to_23,	ready_23_to_22;
wire    [`DW-1:0]   data_23_to_24,	data_24_to_23;
wire                valid_23_to_24,	valid_24_to_23;
wire                ready_23_to_24,	ready_24_to_23;
wire    [`DW-1:0]   data_24_to_25,	data_25_to_24;
wire                valid_24_to_25,	valid_25_to_24;
wire                ready_24_to_25,	ready_25_to_24;
wire    [`DW-1:0]   data_25_to_26,	data_26_to_25;
wire                valid_25_to_26,	valid_26_to_25;
wire                ready_25_to_26,	ready_26_to_25;
wire    [`DW-1:0]   data_26_to_27,	data_27_to_26;
wire                valid_26_to_27,	valid_27_to_26;
wire                ready_26_to_27,	ready_27_to_26;
wire    [`DW-1:0]   data_27_to_28,	data_28_to_27;
wire                valid_27_to_28,	valid_28_to_27;
wire                ready_27_to_28,	ready_28_to_27;
wire    [`DW-1:0]   data_28_to_29,	data_29_to_28;
wire                valid_28_to_29,	valid_29_to_28;
wire                ready_28_to_29,	ready_29_to_28;
wire    [`DW-1:0]   data_30_to_31,	data_31_to_30;
wire                valid_30_to_31,	valid_31_to_30;
wire                ready_30_to_31,	ready_31_to_30;
wire    [`DW-1:0]   data_31_to_32,	data_32_to_31;
wire                valid_31_to_32,	valid_32_to_31;
wire                ready_31_to_32,	ready_32_to_31;
wire    [`DW-1:0]   data_32_to_33,	data_33_to_32;
wire                valid_32_to_33,	valid_33_to_32;
wire                ready_32_to_33,	ready_33_to_32;
wire    [`DW-1:0]   data_33_to_34,	data_34_to_33;
wire                valid_33_to_34,	valid_34_to_33;
wire                ready_33_to_34,	ready_34_to_33;
wire    [`DW-1:0]   data_34_to_35,	data_35_to_34;
wire                valid_34_to_35,	valid_35_to_34;
wire                ready_34_to_35,	ready_35_to_34;
wire    [`DW-1:0]   data_35_to_36,	data_36_to_35;
wire                valid_35_to_36,	valid_36_to_35;
wire                ready_35_to_36,	ready_36_to_35;
wire    [`DW-1:0]   data_36_to_37,	data_37_to_36;
wire                valid_36_to_37,	valid_37_to_36;
wire                ready_36_to_37,	ready_37_to_36;
wire    [`DW-1:0]   data_37_to_38,	data_38_to_37;
wire                valid_37_to_38,	valid_38_to_37;
wire                ready_37_to_38,	ready_38_to_37;
wire    [`DW-1:0]   data_38_to_39,	data_39_to_38;
wire                valid_38_to_39,	valid_39_to_38;
wire                ready_38_to_39,	ready_39_to_38;
wire    [`DW-1:0]   data_40_to_41,	data_41_to_40;
wire                valid_40_to_41,	valid_41_to_40;
wire                ready_40_to_41,	ready_41_to_40;
wire    [`DW-1:0]   data_41_to_42,	data_42_to_41;
wire                valid_41_to_42,	valid_42_to_41;
wire                ready_41_to_42,	ready_42_to_41;
wire    [`DW-1:0]   data_42_to_43,	data_43_to_42;
wire                valid_42_to_43,	valid_43_to_42;
wire                ready_42_to_43,	ready_43_to_42;
wire    [`DW-1:0]   data_43_to_44,	data_44_to_43;
wire                valid_43_to_44,	valid_44_to_43;
wire                ready_43_to_44,	ready_44_to_43;
wire    [`DW-1:0]   data_44_to_45,	data_45_to_44;
wire                valid_44_to_45,	valid_45_to_44;
wire                ready_44_to_45,	ready_45_to_44;
wire    [`DW-1:0]   data_45_to_46,	data_46_to_45;
wire                valid_45_to_46,	valid_46_to_45;
wire                ready_45_to_46,	ready_46_to_45;
wire    [`DW-1:0]   data_46_to_47,	data_47_to_46;
wire                valid_46_to_47,	valid_47_to_46;
wire                ready_46_to_47,	ready_47_to_46;
wire    [`DW-1:0]   data_47_to_48,	data_48_to_47;
wire                valid_47_to_48,	valid_48_to_47;
wire                ready_47_to_48,	ready_48_to_47;
wire    [`DW-1:0]   data_48_to_49,	data_49_to_48;
wire                valid_48_to_49,	valid_49_to_48;
wire                ready_48_to_49,	ready_49_to_48;
wire    [`DW-1:0]   data_50_to_51,	data_51_to_50;
wire                valid_50_to_51,	valid_51_to_50;
wire                ready_50_to_51,	ready_51_to_50;
wire    [`DW-1:0]   data_51_to_52,	data_52_to_51;
wire                valid_51_to_52,	valid_52_to_51;
wire                ready_51_to_52,	ready_52_to_51;
wire    [`DW-1:0]   data_52_to_53,	data_53_to_52;
wire                valid_52_to_53,	valid_53_to_52;
wire                ready_52_to_53,	ready_53_to_52;
wire    [`DW-1:0]   data_53_to_54,	data_54_to_53;
wire                valid_53_to_54,	valid_54_to_53;
wire                ready_53_to_54,	ready_54_to_53;
wire    [`DW-1:0]   data_54_to_55,	data_55_to_54;
wire                valid_54_to_55,	valid_55_to_54;
wire                ready_54_to_55,	ready_55_to_54;
wire    [`DW-1:0]   data_55_to_56,	data_56_to_55;
wire                valid_55_to_56,	valid_56_to_55;
wire                ready_55_to_56,	ready_56_to_55;
wire    [`DW-1:0]   data_56_to_57,	data_57_to_56;
wire                valid_56_to_57,	valid_57_to_56;
wire                ready_56_to_57,	ready_57_to_56;
wire    [`DW-1:0]   data_57_to_58,	data_58_to_57;
wire                valid_57_to_58,	valid_58_to_57;
wire                ready_57_to_58,	ready_58_to_57;
wire    [`DW-1:0]   data_58_to_59,	data_59_to_58;
wire                valid_58_to_59,	valid_59_to_58;
wire                ready_58_to_59,	ready_59_to_58;
wire    [`DW-1:0]   data_60_to_61,	data_61_to_60;
wire                valid_60_to_61,	valid_61_to_60;
wire                ready_60_to_61,	ready_61_to_60;
wire    [`DW-1:0]   data_61_to_62,	data_62_to_61;
wire                valid_61_to_62,	valid_62_to_61;
wire                ready_61_to_62,	ready_62_to_61;
wire    [`DW-1:0]   data_62_to_63,	data_63_to_62;
wire                valid_62_to_63,	valid_63_to_62;
wire                ready_62_to_63,	ready_63_to_62;
wire    [`DW-1:0]   data_63_to_64,	data_64_to_63;
wire                valid_63_to_64,	valid_64_to_63;
wire                ready_63_to_64,	ready_64_to_63;
wire    [`DW-1:0]   data_64_to_65,	data_65_to_64;
wire                valid_64_to_65,	valid_65_to_64;
wire                ready_64_to_65,	ready_65_to_64;
wire    [`DW-1:0]   data_65_to_66,	data_66_to_65;
wire                valid_65_to_66,	valid_66_to_65;
wire                ready_65_to_66,	ready_66_to_65;
wire    [`DW-1:0]   data_66_to_67,	data_67_to_66;
wire                valid_66_to_67,	valid_67_to_66;
wire                ready_66_to_67,	ready_67_to_66;
wire    [`DW-1:0]   data_67_to_68,	data_68_to_67;
wire                valid_67_to_68,	valid_68_to_67;
wire                ready_67_to_68,	ready_68_to_67;
wire    [`DW-1:0]   data_68_to_69,	data_69_to_68;
wire                valid_68_to_69,	valid_69_to_68;
wire                ready_68_to_69,	ready_69_to_68;
wire    [`DW-1:0]   data_70_to_71,	data_71_to_70;
wire                valid_70_to_71,	valid_71_to_70;
wire                ready_70_to_71,	ready_71_to_70;
wire    [`DW-1:0]   data_71_to_72,	data_72_to_71;
wire                valid_71_to_72,	valid_72_to_71;
wire                ready_71_to_72,	ready_72_to_71;
wire    [`DW-1:0]   data_72_to_73,	data_73_to_72;
wire                valid_72_to_73,	valid_73_to_72;
wire                ready_72_to_73,	ready_73_to_72;
wire    [`DW-1:0]   data_73_to_74,	data_74_to_73;
wire                valid_73_to_74,	valid_74_to_73;
wire                ready_73_to_74,	ready_74_to_73;
wire    [`DW-1:0]   data_74_to_75,	data_75_to_74;
wire                valid_74_to_75,	valid_75_to_74;
wire                ready_74_to_75,	ready_75_to_74;
wire    [`DW-1:0]   data_75_to_76,	data_76_to_75;
wire                valid_75_to_76,	valid_76_to_75;
wire                ready_75_to_76,	ready_76_to_75;
wire    [`DW-1:0]   data_76_to_77,	data_77_to_76;
wire                valid_76_to_77,	valid_77_to_76;
wire                ready_76_to_77,	ready_77_to_76;
wire    [`DW-1:0]   data_77_to_78,	data_78_to_77;
wire                valid_77_to_78,	valid_78_to_77;
wire                ready_77_to_78,	ready_78_to_77;
wire    [`DW-1:0]   data_78_to_79,	data_79_to_78;
wire                valid_78_to_79,	valid_79_to_78;
wire                ready_78_to_79,	ready_79_to_78;
wire    [`DW-1:0]   data_80_to_81,	data_81_to_80;
wire                valid_80_to_81,	valid_81_to_80;
wire                ready_80_to_81,	ready_81_to_80;
wire    [`DW-1:0]   data_81_to_82,	data_82_to_81;
wire                valid_81_to_82,	valid_82_to_81;
wire                ready_81_to_82,	ready_82_to_81;
wire    [`DW-1:0]   data_82_to_83,	data_83_to_82;
wire                valid_82_to_83,	valid_83_to_82;
wire                ready_82_to_83,	ready_83_to_82;
wire    [`DW-1:0]   data_83_to_84,	data_84_to_83;
wire                valid_83_to_84,	valid_84_to_83;
wire                ready_83_to_84,	ready_84_to_83;
wire    [`DW-1:0]   data_84_to_85,	data_85_to_84;
wire                valid_84_to_85,	valid_85_to_84;
wire                ready_84_to_85,	ready_85_to_84;
wire    [`DW-1:0]   data_85_to_86,	data_86_to_85;
wire                valid_85_to_86,	valid_86_to_85;
wire                ready_85_to_86,	ready_86_to_85;
wire    [`DW-1:0]   data_86_to_87,	data_87_to_86;
wire                valid_86_to_87,	valid_87_to_86;
wire                ready_86_to_87,	ready_87_to_86;
wire    [`DW-1:0]   data_87_to_88,	data_88_to_87;
wire                valid_87_to_88,	valid_88_to_87;
wire                ready_87_to_88,	ready_88_to_87;
wire    [`DW-1:0]   data_88_to_89,	data_89_to_88;
wire                valid_88_to_89,	valid_89_to_88;
wire                ready_88_to_89,	ready_89_to_88;
wire    [`DW-1:0]   data_90_to_91,	data_91_to_90;
wire                valid_90_to_91,	valid_91_to_90;
wire                ready_90_to_91,	ready_91_to_90;
wire    [`DW-1:0]   data_91_to_92,	data_92_to_91;
wire                valid_91_to_92,	valid_92_to_91;
wire                ready_91_to_92,	ready_92_to_91;
wire    [`DW-1:0]   data_92_to_93,	data_93_to_92;
wire                valid_92_to_93,	valid_93_to_92;
wire                ready_92_to_93,	ready_93_to_92;
wire    [`DW-1:0]   data_93_to_94,	data_94_to_93;
wire                valid_93_to_94,	valid_94_to_93;
wire                ready_93_to_94,	ready_94_to_93;
wire    [`DW-1:0]   data_94_to_95,	data_95_to_94;
wire                valid_94_to_95,	valid_95_to_94;
wire                ready_94_to_95,	ready_95_to_94;
wire    [`DW-1:0]   data_95_to_96,	data_96_to_95;
wire                valid_95_to_96,	valid_96_to_95;
wire                ready_95_to_96,	ready_96_to_95;
wire    [`DW-1:0]   data_96_to_97,	data_97_to_96;
wire                valid_96_to_97,	valid_97_to_96;
wire                ready_96_to_97,	ready_97_to_96;
wire    [`DW-1:0]   data_97_to_98,	data_98_to_97;
wire                valid_97_to_98,	valid_98_to_97;
wire                ready_97_to_98,	ready_98_to_97;
wire    [`DW-1:0]   data_98_to_99,	data_99_to_98;
wire                valid_98_to_99,	valid_99_to_98;
wire                ready_98_to_99,	ready_99_to_98;
wire    [`DW-1:0]   data_100_to_101,	data_101_to_100;
wire                valid_100_to_101,	valid_101_to_100;
wire                ready_100_to_101,	ready_101_to_100;
wire    [`DW-1:0]   data_101_to_102,	data_102_to_101;
wire                valid_101_to_102,	valid_102_to_101;
wire                ready_101_to_102,	ready_102_to_101;
wire    [`DW-1:0]   data_102_to_103,	data_103_to_102;
wire                valid_102_to_103,	valid_103_to_102;
wire                ready_102_to_103,	ready_103_to_102;
wire    [`DW-1:0]   data_103_to_104,	data_104_to_103;
wire                valid_103_to_104,	valid_104_to_103;
wire                ready_103_to_104,	ready_104_to_103;
wire    [`DW-1:0]   data_104_to_105,	data_105_to_104;
wire                valid_104_to_105,	valid_105_to_104;
wire                ready_104_to_105,	ready_105_to_104;
wire    [`DW-1:0]   data_105_to_106,	data_106_to_105;
wire                valid_105_to_106,	valid_106_to_105;
wire                ready_105_to_106,	ready_106_to_105;
wire    [`DW-1:0]   data_106_to_107,	data_107_to_106;
wire                valid_106_to_107,	valid_107_to_106;
wire                ready_106_to_107,	ready_107_to_106;
wire    [`DW-1:0]   data_107_to_108,	data_108_to_107;
wire                valid_107_to_108,	valid_108_to_107;
wire                ready_107_to_108,	ready_108_to_107;
wire    [`DW-1:0]   data_108_to_109,	data_109_to_108;
wire                valid_108_to_109,	valid_109_to_108;
wire                ready_108_to_109,	ready_109_to_108;
wire    [`DW-1:0]   data_110_to_111,	data_111_to_110;
wire                valid_110_to_111,	valid_111_to_110;
wire                ready_110_to_111,	ready_111_to_110;
wire    [`DW-1:0]   data_111_to_112,	data_112_to_111;
wire                valid_111_to_112,	valid_112_to_111;
wire                ready_111_to_112,	ready_112_to_111;
wire    [`DW-1:0]   data_112_to_113,	data_113_to_112;
wire                valid_112_to_113,	valid_113_to_112;
wire                ready_112_to_113,	ready_113_to_112;
wire    [`DW-1:0]   data_113_to_114,	data_114_to_113;
wire                valid_113_to_114,	valid_114_to_113;
wire                ready_113_to_114,	ready_114_to_113;
wire    [`DW-1:0]   data_114_to_115,	data_115_to_114;
wire                valid_114_to_115,	valid_115_to_114;
wire                ready_114_to_115,	ready_115_to_114;
wire    [`DW-1:0]   data_115_to_116,	data_116_to_115;
wire                valid_115_to_116,	valid_116_to_115;
wire                ready_115_to_116,	ready_116_to_115;
wire    [`DW-1:0]   data_116_to_117,	data_117_to_116;
wire                valid_116_to_117,	valid_117_to_116;
wire                ready_116_to_117,	ready_117_to_116;
wire    [`DW-1:0]   data_117_to_118,	data_118_to_117;
wire                valid_117_to_118,	valid_118_to_117;
wire                ready_117_to_118,	ready_118_to_117;
wire    [`DW-1:0]   data_118_to_119,	data_119_to_118;
wire                valid_118_to_119,	valid_119_to_118;
wire                ready_118_to_119,	ready_119_to_118;
wire    [`DW-1:0]   data_120_to_121,	data_121_to_120;
wire                valid_120_to_121,	valid_121_to_120;
wire                ready_120_to_121,	ready_121_to_120;
wire    [`DW-1:0]   data_121_to_122,	data_122_to_121;
wire                valid_121_to_122,	valid_122_to_121;
wire                ready_121_to_122,	ready_122_to_121;
wire    [`DW-1:0]   data_122_to_123,	data_123_to_122;
wire                valid_122_to_123,	valid_123_to_122;
wire                ready_122_to_123,	ready_123_to_122;
wire    [`DW-1:0]   data_123_to_124,	data_124_to_123;
wire                valid_123_to_124,	valid_124_to_123;
wire                ready_123_to_124,	ready_124_to_123;
wire    [`DW-1:0]   data_124_to_125,	data_125_to_124;
wire                valid_124_to_125,	valid_125_to_124;
wire                ready_124_to_125,	ready_125_to_124;
wire    [`DW-1:0]   data_125_to_126,	data_126_to_125;
wire                valid_125_to_126,	valid_126_to_125;
wire                ready_125_to_126,	ready_126_to_125;
wire    [`DW-1:0]   data_126_to_127,	data_127_to_126;
wire                valid_126_to_127,	valid_127_to_126;
wire                ready_126_to_127,	ready_127_to_126;
wire    [`DW-1:0]   data_127_to_128,	data_128_to_127;
wire                valid_127_to_128,	valid_128_to_127;
wire                ready_127_to_128,	ready_128_to_127;
wire    [`DW-1:0]   data_128_to_129,	data_129_to_128;
wire                valid_128_to_129,	valid_129_to_128;
wire                ready_128_to_129,	ready_129_to_128;
wire    [`DW-1:0]   data_130_to_131,	data_131_to_130;
wire                valid_130_to_131,	valid_131_to_130;
wire                ready_130_to_131,	ready_131_to_130;
wire    [`DW-1:0]   data_131_to_132,	data_132_to_131;
wire                valid_131_to_132,	valid_132_to_131;
wire                ready_131_to_132,	ready_132_to_131;
wire    [`DW-1:0]   data_132_to_133,	data_133_to_132;
wire                valid_132_to_133,	valid_133_to_132;
wire                ready_132_to_133,	ready_133_to_132;
wire    [`DW-1:0]   data_133_to_134,	data_134_to_133;
wire                valid_133_to_134,	valid_134_to_133;
wire                ready_133_to_134,	ready_134_to_133;
wire    [`DW-1:0]   data_134_to_135,	data_135_to_134;
wire                valid_134_to_135,	valid_135_to_134;
wire                ready_134_to_135,	ready_135_to_134;
wire    [`DW-1:0]   data_135_to_136,	data_136_to_135;
wire                valid_135_to_136,	valid_136_to_135;
wire                ready_135_to_136,	ready_136_to_135;
wire    [`DW-1:0]   data_136_to_137,	data_137_to_136;
wire                valid_136_to_137,	valid_137_to_136;
wire                ready_136_to_137,	ready_137_to_136;
wire    [`DW-1:0]   data_137_to_138,	data_138_to_137;
wire                valid_137_to_138,	valid_138_to_137;
wire                ready_137_to_138,	ready_138_to_137;
wire    [`DW-1:0]   data_138_to_139,	data_139_to_138;
wire                valid_138_to_139,	valid_139_to_138;
wire                ready_138_to_139,	ready_139_to_138;
wire    [`DW-1:0]   data_140_to_141,	data_141_to_140;
wire                valid_140_to_141,	valid_141_to_140;
wire                ready_140_to_141,	ready_141_to_140;
wire    [`DW-1:0]   data_141_to_142,	data_142_to_141;
wire                valid_141_to_142,	valid_142_to_141;
wire                ready_141_to_142,	ready_142_to_141;
wire    [`DW-1:0]   data_142_to_143,	data_143_to_142;
wire                valid_142_to_143,	valid_143_to_142;
wire                ready_142_to_143,	ready_143_to_142;
wire    [`DW-1:0]   data_143_to_144,	data_144_to_143;
wire                valid_143_to_144,	valid_144_to_143;
wire                ready_143_to_144,	ready_144_to_143;
wire    [`DW-1:0]   data_144_to_145,	data_145_to_144;
wire                valid_144_to_145,	valid_145_to_144;
wire                ready_144_to_145,	ready_145_to_144;
wire    [`DW-1:0]   data_145_to_146,	data_146_to_145;
wire                valid_145_to_146,	valid_146_to_145;
wire                ready_145_to_146,	ready_146_to_145;
wire    [`DW-1:0]   data_146_to_147,	data_147_to_146;
wire                valid_146_to_147,	valid_147_to_146;
wire                ready_146_to_147,	ready_147_to_146;
wire    [`DW-1:0]   data_147_to_148,	data_148_to_147;
wire                valid_147_to_148,	valid_148_to_147;
wire                ready_147_to_148,	ready_148_to_147;
wire    [`DW-1:0]   data_148_to_149,	data_149_to_148;
wire                valid_148_to_149,	valid_149_to_148;
wire                ready_148_to_149,	ready_149_to_148;
wire    [`DW-1:0]   data_150_to_151,	data_151_to_150;
wire                valid_150_to_151,	valid_151_to_150;
wire                ready_150_to_151,	ready_151_to_150;
wire    [`DW-1:0]   data_151_to_152,	data_152_to_151;
wire                valid_151_to_152,	valid_152_to_151;
wire                ready_151_to_152,	ready_152_to_151;
wire    [`DW-1:0]   data_152_to_153,	data_153_to_152;
wire                valid_152_to_153,	valid_153_to_152;
wire                ready_152_to_153,	ready_153_to_152;
wire    [`DW-1:0]   data_153_to_154,	data_154_to_153;
wire                valid_153_to_154,	valid_154_to_153;
wire                ready_153_to_154,	ready_154_to_153;
wire    [`DW-1:0]   data_154_to_155,	data_155_to_154;
wire                valid_154_to_155,	valid_155_to_154;
wire                ready_154_to_155,	ready_155_to_154;
wire    [`DW-1:0]   data_155_to_156,	data_156_to_155;
wire                valid_155_to_156,	valid_156_to_155;
wire                ready_155_to_156,	ready_156_to_155;
wire    [`DW-1:0]   data_156_to_157,	data_157_to_156;
wire                valid_156_to_157,	valid_157_to_156;
wire                ready_156_to_157,	ready_157_to_156;
wire    [`DW-1:0]   data_157_to_158,	data_158_to_157;
wire                valid_157_to_158,	valid_158_to_157;
wire                ready_157_to_158,	ready_158_to_157;
wire    [`DW-1:0]   data_158_to_159,	data_159_to_158;
wire                valid_158_to_159,	valid_159_to_158;
wire                ready_158_to_159,	ready_159_to_158;
wire    [`DW-1:0]   data_160_to_161,	data_161_to_160;
wire                valid_160_to_161,	valid_161_to_160;
wire                ready_160_to_161,	ready_161_to_160;
wire    [`DW-1:0]   data_161_to_162,	data_162_to_161;
wire                valid_161_to_162,	valid_162_to_161;
wire                ready_161_to_162,	ready_162_to_161;
wire    [`DW-1:0]   data_162_to_163,	data_163_to_162;
wire                valid_162_to_163,	valid_163_to_162;
wire                ready_162_to_163,	ready_163_to_162;
wire    [`DW-1:0]   data_163_to_164,	data_164_to_163;
wire                valid_163_to_164,	valid_164_to_163;
wire                ready_163_to_164,	ready_164_to_163;
wire    [`DW-1:0]   data_164_to_165,	data_165_to_164;
wire                valid_164_to_165,	valid_165_to_164;
wire                ready_164_to_165,	ready_165_to_164;
wire    [`DW-1:0]   data_165_to_166,	data_166_to_165;
wire                valid_165_to_166,	valid_166_to_165;
wire                ready_165_to_166,	ready_166_to_165;
wire    [`DW-1:0]   data_166_to_167,	data_167_to_166;
wire                valid_166_to_167,	valid_167_to_166;
wire                ready_166_to_167,	ready_167_to_166;
wire    [`DW-1:0]   data_167_to_168,	data_168_to_167;
wire                valid_167_to_168,	valid_168_to_167;
wire                ready_167_to_168,	ready_168_to_167;
wire    [`DW-1:0]   data_168_to_169,	data_169_to_168;
wire                valid_168_to_169,	valid_169_to_168;
wire                ready_168_to_169,	ready_169_to_168;
wire    [`DW-1:0]   data_170_to_171,	data_171_to_170;
wire                valid_170_to_171,	valid_171_to_170;
wire                ready_170_to_171,	ready_171_to_170;
wire    [`DW-1:0]   data_171_to_172,	data_172_to_171;
wire                valid_171_to_172,	valid_172_to_171;
wire                ready_171_to_172,	ready_172_to_171;
wire    [`DW-1:0]   data_172_to_173,	data_173_to_172;
wire                valid_172_to_173,	valid_173_to_172;
wire                ready_172_to_173,	ready_173_to_172;
wire    [`DW-1:0]   data_173_to_174,	data_174_to_173;
wire                valid_173_to_174,	valid_174_to_173;
wire                ready_173_to_174,	ready_174_to_173;
wire    [`DW-1:0]   data_174_to_175,	data_175_to_174;
wire                valid_174_to_175,	valid_175_to_174;
wire                ready_174_to_175,	ready_175_to_174;
wire    [`DW-1:0]   data_175_to_176,	data_176_to_175;
wire                valid_175_to_176,	valid_176_to_175;
wire                ready_175_to_176,	ready_176_to_175;
wire    [`DW-1:0]   data_176_to_177,	data_177_to_176;
wire                valid_176_to_177,	valid_177_to_176;
wire                ready_176_to_177,	ready_177_to_176;
wire    [`DW-1:0]   data_177_to_178,	data_178_to_177;
wire                valid_177_to_178,	valid_178_to_177;
wire                ready_177_to_178,	ready_178_to_177;
wire    [`DW-1:0]   data_178_to_179,	data_179_to_178;
wire                valid_178_to_179,	valid_179_to_178;
wire                ready_178_to_179,	ready_179_to_178;
wire    [`DW-1:0]   data_180_to_181,	data_181_to_180;
wire                valid_180_to_181,	valid_181_to_180;
wire                ready_180_to_181,	ready_181_to_180;
wire    [`DW-1:0]   data_181_to_182,	data_182_to_181;
wire                valid_181_to_182,	valid_182_to_181;
wire                ready_181_to_182,	ready_182_to_181;
wire    [`DW-1:0]   data_182_to_183,	data_183_to_182;
wire                valid_182_to_183,	valid_183_to_182;
wire                ready_182_to_183,	ready_183_to_182;
wire    [`DW-1:0]   data_183_to_184,	data_184_to_183;
wire                valid_183_to_184,	valid_184_to_183;
wire                ready_183_to_184,	ready_184_to_183;
wire    [`DW-1:0]   data_184_to_185,	data_185_to_184;
wire                valid_184_to_185,	valid_185_to_184;
wire                ready_184_to_185,	ready_185_to_184;
wire    [`DW-1:0]   data_185_to_186,	data_186_to_185;
wire                valid_185_to_186,	valid_186_to_185;
wire                ready_185_to_186,	ready_186_to_185;
wire    [`DW-1:0]   data_186_to_187,	data_187_to_186;
wire                valid_186_to_187,	valid_187_to_186;
wire                ready_186_to_187,	ready_187_to_186;
wire    [`DW-1:0]   data_187_to_188,	data_188_to_187;
wire                valid_187_to_188,	valid_188_to_187;
wire                ready_187_to_188,	ready_188_to_187;
wire    [`DW-1:0]   data_188_to_189,	data_189_to_188;
wire                valid_188_to_189,	valid_189_to_188;
wire                ready_188_to_189,	ready_189_to_188;
wire    [`DW-1:0]   data_190_to_191,	data_191_to_190;
wire                valid_190_to_191,	valid_191_to_190;
wire                ready_190_to_191,	ready_191_to_190;
wire    [`DW-1:0]   data_191_to_192,	data_192_to_191;
wire                valid_191_to_192,	valid_192_to_191;
wire                ready_191_to_192,	ready_192_to_191;
wire    [`DW-1:0]   data_192_to_193,	data_193_to_192;
wire                valid_192_to_193,	valid_193_to_192;
wire                ready_192_to_193,	ready_193_to_192;
wire    [`DW-1:0]   data_193_to_194,	data_194_to_193;
wire                valid_193_to_194,	valid_194_to_193;
wire                ready_193_to_194,	ready_194_to_193;
wire    [`DW-1:0]   data_194_to_195,	data_195_to_194;
wire                valid_194_to_195,	valid_195_to_194;
wire                ready_194_to_195,	ready_195_to_194;
wire    [`DW-1:0]   data_195_to_196,	data_196_to_195;
wire                valid_195_to_196,	valid_196_to_195;
wire                ready_195_to_196,	ready_196_to_195;
wire    [`DW-1:0]   data_196_to_197,	data_197_to_196;
wire                valid_196_to_197,	valid_197_to_196;
wire                ready_196_to_197,	ready_197_to_196;
wire    [`DW-1:0]   data_197_to_198,	data_198_to_197;
wire                valid_197_to_198,	valid_198_to_197;
wire                ready_197_to_198,	ready_198_to_197;
wire    [`DW-1:0]   data_198_to_199,	data_199_to_198;
wire                valid_198_to_199,	valid_199_to_198;
wire                ready_198_to_199,	ready_199_to_198;
wire    [`DW-1:0]   data_200_to_201,	data_201_to_200;
wire                valid_200_to_201,	valid_201_to_200;
wire                ready_200_to_201,	ready_201_to_200;
wire    [`DW-1:0]   data_201_to_202,	data_202_to_201;
wire                valid_201_to_202,	valid_202_to_201;
wire                ready_201_to_202,	ready_202_to_201;
wire    [`DW-1:0]   data_202_to_203,	data_203_to_202;
wire                valid_202_to_203,	valid_203_to_202;
wire                ready_202_to_203,	ready_203_to_202;
wire    [`DW-1:0]   data_203_to_204,	data_204_to_203;
wire                valid_203_to_204,	valid_204_to_203;
wire                ready_203_to_204,	ready_204_to_203;
wire    [`DW-1:0]   data_204_to_205,	data_205_to_204;
wire                valid_204_to_205,	valid_205_to_204;
wire                ready_204_to_205,	ready_205_to_204;
wire    [`DW-1:0]   data_205_to_206,	data_206_to_205;
wire                valid_205_to_206,	valid_206_to_205;
wire                ready_205_to_206,	ready_206_to_205;
wire    [`DW-1:0]   data_206_to_207,	data_207_to_206;
wire                valid_206_to_207,	valid_207_to_206;
wire                ready_206_to_207,	ready_207_to_206;
wire    [`DW-1:0]   data_207_to_208,	data_208_to_207;
wire                valid_207_to_208,	valid_208_to_207;
wire                ready_207_to_208,	ready_208_to_207;
wire    [`DW-1:0]   data_208_to_209,	data_209_to_208;
wire                valid_208_to_209,	valid_209_to_208;
wire                ready_208_to_209,	ready_209_to_208;
wire    [`DW-1:0]   data_210_to_211,	data_211_to_210;
wire                valid_210_to_211,	valid_211_to_210;
wire                ready_210_to_211,	ready_211_to_210;
wire    [`DW-1:0]   data_211_to_212,	data_212_to_211;
wire                valid_211_to_212,	valid_212_to_211;
wire                ready_211_to_212,	ready_212_to_211;
wire    [`DW-1:0]   data_212_to_213,	data_213_to_212;
wire                valid_212_to_213,	valid_213_to_212;
wire                ready_212_to_213,	ready_213_to_212;
wire    [`DW-1:0]   data_213_to_214,	data_214_to_213;
wire                valid_213_to_214,	valid_214_to_213;
wire                ready_213_to_214,	ready_214_to_213;
wire    [`DW-1:0]   data_214_to_215,	data_215_to_214;
wire                valid_214_to_215,	valid_215_to_214;
wire                ready_214_to_215,	ready_215_to_214;
wire    [`DW-1:0]   data_215_to_216,	data_216_to_215;
wire                valid_215_to_216,	valid_216_to_215;
wire                ready_215_to_216,	ready_216_to_215;
wire    [`DW-1:0]   data_216_to_217,	data_217_to_216;
wire                valid_216_to_217,	valid_217_to_216;
wire                ready_216_to_217,	ready_217_to_216;
wire    [`DW-1:0]   data_217_to_218,	data_218_to_217;
wire                valid_217_to_218,	valid_218_to_217;
wire                ready_217_to_218,	ready_218_to_217;
wire    [`DW-1:0]   data_218_to_219,	data_219_to_218;
wire                valid_218_to_219,	valid_219_to_218;
wire                ready_218_to_219,	ready_219_to_218;
wire    [`DW-1:0]   data_220_to_221,	data_221_to_220;
wire                valid_220_to_221,	valid_221_to_220;
wire                ready_220_to_221,	ready_221_to_220;
wire    [`DW-1:0]   data_221_to_222,	data_222_to_221;
wire                valid_221_to_222,	valid_222_to_221;
wire                ready_221_to_222,	ready_222_to_221;
wire    [`DW-1:0]   data_222_to_223,	data_223_to_222;
wire                valid_222_to_223,	valid_223_to_222;
wire                ready_222_to_223,	ready_223_to_222;
wire    [`DW-1:0]   data_223_to_224,	data_224_to_223;
wire                valid_223_to_224,	valid_224_to_223;
wire                ready_223_to_224,	ready_224_to_223;
wire    [`DW-1:0]   data_224_to_225,	data_225_to_224;
wire                valid_224_to_225,	valid_225_to_224;
wire                ready_224_to_225,	ready_225_to_224;
wire    [`DW-1:0]   data_225_to_226,	data_226_to_225;
wire                valid_225_to_226,	valid_226_to_225;
wire                ready_225_to_226,	ready_226_to_225;
wire    [`DW-1:0]   data_226_to_227,	data_227_to_226;
wire                valid_226_to_227,	valid_227_to_226;
wire                ready_226_to_227,	ready_227_to_226;
wire    [`DW-1:0]   data_227_to_228,	data_228_to_227;
wire                valid_227_to_228,	valid_228_to_227;
wire                ready_227_to_228,	ready_228_to_227;
wire    [`DW-1:0]   data_228_to_229,	data_229_to_228;
wire                valid_228_to_229,	valid_229_to_228;
wire                ready_228_to_229,	ready_229_to_228;
wire    [`DW-1:0]   data_230_to_231,	data_231_to_230;
wire                valid_230_to_231,	valid_231_to_230;
wire                ready_230_to_231,	ready_231_to_230;
wire    [`DW-1:0]   data_231_to_232,	data_232_to_231;
wire                valid_231_to_232,	valid_232_to_231;
wire                ready_231_to_232,	ready_232_to_231;
wire    [`DW-1:0]   data_232_to_233,	data_233_to_232;
wire                valid_232_to_233,	valid_233_to_232;
wire                ready_232_to_233,	ready_233_to_232;
wire    [`DW-1:0]   data_233_to_234,	data_234_to_233;
wire                valid_233_to_234,	valid_234_to_233;
wire                ready_233_to_234,	ready_234_to_233;
wire    [`DW-1:0]   data_234_to_235,	data_235_to_234;
wire                valid_234_to_235,	valid_235_to_234;
wire                ready_234_to_235,	ready_235_to_234;
wire    [`DW-1:0]   data_235_to_236,	data_236_to_235;
wire                valid_235_to_236,	valid_236_to_235;
wire                ready_235_to_236,	ready_236_to_235;
wire    [`DW-1:0]   data_236_to_237,	data_237_to_236;
wire                valid_236_to_237,	valid_237_to_236;
wire                ready_236_to_237,	ready_237_to_236;
wire    [`DW-1:0]   data_237_to_238,	data_238_to_237;
wire                valid_237_to_238,	valid_238_to_237;
wire                ready_237_to_238,	ready_238_to_237;
wire    [`DW-1:0]   data_238_to_239,	data_239_to_238;
wire                valid_238_to_239,	valid_239_to_238;
wire                ready_238_to_239,	ready_239_to_238;
wire    [`DW-1:0]   data_240_to_241,	data_241_to_240;
wire                valid_240_to_241,	valid_241_to_240;
wire                ready_240_to_241,	ready_241_to_240;
wire    [`DW-1:0]   data_241_to_242,	data_242_to_241;
wire                valid_241_to_242,	valid_242_to_241;
wire                ready_241_to_242,	ready_242_to_241;
wire    [`DW-1:0]   data_242_to_243,	data_243_to_242;
wire                valid_242_to_243,	valid_243_to_242;
wire                ready_242_to_243,	ready_243_to_242;
wire    [`DW-1:0]   data_243_to_244,	data_244_to_243;
wire                valid_243_to_244,	valid_244_to_243;
wire                ready_243_to_244,	ready_244_to_243;
wire    [`DW-1:0]   data_244_to_245,	data_245_to_244;
wire                valid_244_to_245,	valid_245_to_244;
wire                ready_244_to_245,	ready_245_to_244;
wire    [`DW-1:0]   data_245_to_246,	data_246_to_245;
wire                valid_245_to_246,	valid_246_to_245;
wire                ready_245_to_246,	ready_246_to_245;
wire    [`DW-1:0]   data_246_to_247,	data_247_to_246;
wire                valid_246_to_247,	valid_247_to_246;
wire                ready_246_to_247,	ready_247_to_246;
wire    [`DW-1:0]   data_247_to_248,	data_248_to_247;
wire                valid_247_to_248,	valid_248_to_247;
wire                ready_247_to_248,	ready_248_to_247;
wire    [`DW-1:0]   data_248_to_249,	data_249_to_248;
wire                valid_248_to_249,	valid_249_to_248;
wire                ready_248_to_249,	ready_249_to_248;

//vertical signals
wire    [`DW-1:0]   data_0_to_10_v0,	data_0_to_10_v1;
wire                valid_0_to_10_v0,	valid_0_to_10_v1;
wire                ready_10_to_0_v0,	ready_10_to_0_v1;
wire    [`DW-1:0]   data_10_to_20_v0,	data_10_to_20_v1;
wire                valid_10_to_20_v0,	valid_10_to_20_v1;
wire                ready_20_to_10_v0,	ready_20_to_10_v1;
wire    [`DW-1:0]   data_20_to_30_v0,	data_20_to_30_v1;
wire                valid_20_to_30_v0,	valid_20_to_30_v1;
wire                ready_30_to_20_v0,	ready_30_to_20_v1;
wire    [`DW-1:0]   data_30_to_40_v0,	data_30_to_40_v1;
wire                valid_30_to_40_v0,	valid_30_to_40_v1;
wire                ready_40_to_30_v0,	ready_40_to_30_v1;
wire    [`DW-1:0]   data_40_to_50_v0,	data_40_to_50_v1;
wire                valid_40_to_50_v0,	valid_40_to_50_v1;
wire                ready_50_to_40_v0,	ready_50_to_40_v1;
wire    [`DW-1:0]   data_50_to_60_v0,	data_50_to_60_v1;
wire                valid_50_to_60_v0,	valid_50_to_60_v1;
wire                ready_60_to_50_v0,	ready_60_to_50_v1;
wire    [`DW-1:0]   data_60_to_70_v0,	data_60_to_70_v1;
wire                valid_60_to_70_v0,	valid_60_to_70_v1;
wire                ready_70_to_60_v0,	ready_70_to_60_v1;
wire    [`DW-1:0]   data_70_to_80_v0,	data_70_to_80_v1;
wire                valid_70_to_80_v0,	valid_70_to_80_v1;
wire                ready_80_to_70_v0,	ready_80_to_70_v1;
wire    [`DW-1:0]   data_80_to_90_v0,	data_80_to_90_v1;
wire                valid_80_to_90_v0,	valid_80_to_90_v1;
wire                ready_90_to_80_v0,	ready_90_to_80_v1;
wire    [`DW-1:0]   data_90_to_100_v0,	data_90_to_100_v1;
wire                valid_90_to_100_v0,	valid_90_to_100_v1;
wire                ready_100_to_90_v0,	ready_100_to_90_v1;
wire    [`DW-1:0]   data_100_to_110_v0,	data_100_to_110_v1;
wire                valid_100_to_110_v0,	valid_100_to_110_v1;
wire                ready_110_to_100_v0,	ready_110_to_100_v1;
wire    [`DW-1:0]   data_110_to_120_v0,	data_110_to_120_v1;
wire                valid_110_to_120_v0,	valid_110_to_120_v1;
wire                ready_120_to_110_v0,	ready_120_to_110_v1;
wire    [`DW-1:0]   data_120_to_130_v0,	data_120_to_130_v1;
wire                valid_120_to_130_v0,	valid_120_to_130_v1;
wire                ready_130_to_120_v0,	ready_130_to_120_v1;
wire    [`DW-1:0]   data_130_to_140_v0,	data_130_to_140_v1;
wire                valid_130_to_140_v0,	valid_130_to_140_v1;
wire                ready_140_to_130_v0,	ready_140_to_130_v1;
wire    [`DW-1:0]   data_140_to_150_v0,	data_140_to_150_v1;
wire                valid_140_to_150_v0,	valid_140_to_150_v1;
wire                ready_150_to_140_v0,	ready_150_to_140_v1;
wire    [`DW-1:0]   data_150_to_160_v0,	data_150_to_160_v1;
wire                valid_150_to_160_v0,	valid_150_to_160_v1;
wire                ready_160_to_150_v0,	ready_160_to_150_v1;
wire    [`DW-1:0]   data_160_to_170_v0,	data_160_to_170_v1;
wire                valid_160_to_170_v0,	valid_160_to_170_v1;
wire                ready_170_to_160_v0,	ready_170_to_160_v1;
wire    [`DW-1:0]   data_170_to_180_v0,	data_170_to_180_v1;
wire                valid_170_to_180_v0,	valid_170_to_180_v1;
wire                ready_180_to_170_v0,	ready_180_to_170_v1;
wire    [`DW-1:0]   data_180_to_190_v0,	data_180_to_190_v1;
wire                valid_180_to_190_v0,	valid_180_to_190_v1;
wire                ready_190_to_180_v0,	ready_190_to_180_v1;
wire    [`DW-1:0]   data_190_to_200_v0,	data_190_to_200_v1;
wire                valid_190_to_200_v0,	valid_190_to_200_v1;
wire                ready_200_to_190_v0,	ready_200_to_190_v1;
wire    [`DW-1:0]   data_200_to_210_v0,	data_200_to_210_v1;
wire                valid_200_to_210_v0,	valid_200_to_210_v1;
wire                ready_210_to_200_v0,	ready_210_to_200_v1;
wire    [`DW-1:0]   data_210_to_220_v0,	data_210_to_220_v1;
wire                valid_210_to_220_v0,	valid_210_to_220_v1;
wire                ready_220_to_210_v0,	ready_220_to_210_v1;
wire    [`DW-1:0]   data_220_to_230_v0,	data_220_to_230_v1;
wire                valid_220_to_230_v0,	valid_220_to_230_v1;
wire                ready_230_to_220_v0,	ready_230_to_220_v1;
wire    [`DW-1:0]   data_230_to_240_v0,	data_230_to_240_v1;
wire                valid_230_to_240_v0,	valid_230_to_240_v1;
wire                ready_240_to_230_v0,	ready_240_to_230_v1;
wire    [`DW-1:0]   data_1_to_11_v0,	data_1_to_11_v1;
wire                valid_1_to_11_v0,	valid_1_to_11_v1;
wire                ready_11_to_1_v0,	ready_11_to_1_v1;
wire    [`DW-1:0]   data_11_to_21_v0,	data_11_to_21_v1;
wire                valid_11_to_21_v0,	valid_11_to_21_v1;
wire                ready_21_to_11_v0,	ready_21_to_11_v1;
wire    [`DW-1:0]   data_21_to_31_v0,	data_21_to_31_v1;
wire                valid_21_to_31_v0,	valid_21_to_31_v1;
wire                ready_31_to_21_v0,	ready_31_to_21_v1;
wire    [`DW-1:0]   data_31_to_41_v0,	data_31_to_41_v1;
wire                valid_31_to_41_v0,	valid_31_to_41_v1;
wire                ready_41_to_31_v0,	ready_41_to_31_v1;
wire    [`DW-1:0]   data_41_to_51_v0,	data_41_to_51_v1;
wire                valid_41_to_51_v0,	valid_41_to_51_v1;
wire                ready_51_to_41_v0,	ready_51_to_41_v1;
wire    [`DW-1:0]   data_51_to_61_v0,	data_51_to_61_v1;
wire                valid_51_to_61_v0,	valid_51_to_61_v1;
wire                ready_61_to_51_v0,	ready_61_to_51_v1;
wire    [`DW-1:0]   data_61_to_71_v0,	data_61_to_71_v1;
wire                valid_61_to_71_v0,	valid_61_to_71_v1;
wire                ready_71_to_61_v0,	ready_71_to_61_v1;
wire    [`DW-1:0]   data_71_to_81_v0,	data_71_to_81_v1;
wire                valid_71_to_81_v0,	valid_71_to_81_v1;
wire                ready_81_to_71_v0,	ready_81_to_71_v1;
wire    [`DW-1:0]   data_81_to_91_v0,	data_81_to_91_v1;
wire                valid_81_to_91_v0,	valid_81_to_91_v1;
wire                ready_91_to_81_v0,	ready_91_to_81_v1;
wire    [`DW-1:0]   data_91_to_101_v0,	data_91_to_101_v1;
wire                valid_91_to_101_v0,	valid_91_to_101_v1;
wire                ready_101_to_91_v0,	ready_101_to_91_v1;
wire    [`DW-1:0]   data_101_to_111_v0,	data_101_to_111_v1;
wire                valid_101_to_111_v0,	valid_101_to_111_v1;
wire                ready_111_to_101_v0,	ready_111_to_101_v1;
wire    [`DW-1:0]   data_111_to_121_v0,	data_111_to_121_v1;
wire                valid_111_to_121_v0,	valid_111_to_121_v1;
wire                ready_121_to_111_v0,	ready_121_to_111_v1;
wire    [`DW-1:0]   data_121_to_131_v0,	data_121_to_131_v1;
wire                valid_121_to_131_v0,	valid_121_to_131_v1;
wire                ready_131_to_121_v0,	ready_131_to_121_v1;
wire    [`DW-1:0]   data_131_to_141_v0,	data_131_to_141_v1;
wire                valid_131_to_141_v0,	valid_131_to_141_v1;
wire                ready_141_to_131_v0,	ready_141_to_131_v1;
wire    [`DW-1:0]   data_141_to_151_v0,	data_141_to_151_v1;
wire                valid_141_to_151_v0,	valid_141_to_151_v1;
wire                ready_151_to_141_v0,	ready_151_to_141_v1;
wire    [`DW-1:0]   data_151_to_161_v0,	data_151_to_161_v1;
wire                valid_151_to_161_v0,	valid_151_to_161_v1;
wire                ready_161_to_151_v0,	ready_161_to_151_v1;
wire    [`DW-1:0]   data_161_to_171_v0,	data_161_to_171_v1;
wire                valid_161_to_171_v0,	valid_161_to_171_v1;
wire                ready_171_to_161_v0,	ready_171_to_161_v1;
wire    [`DW-1:0]   data_171_to_181_v0,	data_171_to_181_v1;
wire                valid_171_to_181_v0,	valid_171_to_181_v1;
wire                ready_181_to_171_v0,	ready_181_to_171_v1;
wire    [`DW-1:0]   data_181_to_191_v0,	data_181_to_191_v1;
wire                valid_181_to_191_v0,	valid_181_to_191_v1;
wire                ready_191_to_181_v0,	ready_191_to_181_v1;
wire    [`DW-1:0]   data_191_to_201_v0,	data_191_to_201_v1;
wire                valid_191_to_201_v0,	valid_191_to_201_v1;
wire                ready_201_to_191_v0,	ready_201_to_191_v1;
wire    [`DW-1:0]   data_201_to_211_v0,	data_201_to_211_v1;
wire                valid_201_to_211_v0,	valid_201_to_211_v1;
wire                ready_211_to_201_v0,	ready_211_to_201_v1;
wire    [`DW-1:0]   data_211_to_221_v0,	data_211_to_221_v1;
wire                valid_211_to_221_v0,	valid_211_to_221_v1;
wire                ready_221_to_211_v0,	ready_221_to_211_v1;
wire    [`DW-1:0]   data_221_to_231_v0,	data_221_to_231_v1;
wire                valid_221_to_231_v0,	valid_221_to_231_v1;
wire                ready_231_to_221_v0,	ready_231_to_221_v1;
wire    [`DW-1:0]   data_231_to_241_v0,	data_231_to_241_v1;
wire                valid_231_to_241_v0,	valid_231_to_241_v1;
wire                ready_241_to_231_v0,	ready_241_to_231_v1;
wire    [`DW-1:0]   data_2_to_12_v0,	data_2_to_12_v1;
wire                valid_2_to_12_v0,	valid_2_to_12_v1;
wire                ready_12_to_2_v0,	ready_12_to_2_v1;
wire    [`DW-1:0]   data_12_to_22_v0,	data_12_to_22_v1;
wire                valid_12_to_22_v0,	valid_12_to_22_v1;
wire                ready_22_to_12_v0,	ready_22_to_12_v1;
wire    [`DW-1:0]   data_22_to_32_v0,	data_22_to_32_v1;
wire                valid_22_to_32_v0,	valid_22_to_32_v1;
wire                ready_32_to_22_v0,	ready_32_to_22_v1;
wire    [`DW-1:0]   data_32_to_42_v0,	data_32_to_42_v1;
wire                valid_32_to_42_v0,	valid_32_to_42_v1;
wire                ready_42_to_32_v0,	ready_42_to_32_v1;
wire    [`DW-1:0]   data_42_to_52_v0,	data_42_to_52_v1;
wire                valid_42_to_52_v0,	valid_42_to_52_v1;
wire                ready_52_to_42_v0,	ready_52_to_42_v1;
wire    [`DW-1:0]   data_52_to_62_v0,	data_52_to_62_v1;
wire                valid_52_to_62_v0,	valid_52_to_62_v1;
wire                ready_62_to_52_v0,	ready_62_to_52_v1;
wire    [`DW-1:0]   data_62_to_72_v0,	data_62_to_72_v1;
wire                valid_62_to_72_v0,	valid_62_to_72_v1;
wire                ready_72_to_62_v0,	ready_72_to_62_v1;
wire    [`DW-1:0]   data_72_to_82_v0,	data_72_to_82_v1;
wire                valid_72_to_82_v0,	valid_72_to_82_v1;
wire                ready_82_to_72_v0,	ready_82_to_72_v1;
wire    [`DW-1:0]   data_82_to_92_v0,	data_82_to_92_v1;
wire                valid_82_to_92_v0,	valid_82_to_92_v1;
wire                ready_92_to_82_v0,	ready_92_to_82_v1;
wire    [`DW-1:0]   data_92_to_102_v0,	data_92_to_102_v1;
wire                valid_92_to_102_v0,	valid_92_to_102_v1;
wire                ready_102_to_92_v0,	ready_102_to_92_v1;
wire    [`DW-1:0]   data_102_to_112_v0,	data_102_to_112_v1;
wire                valid_102_to_112_v0,	valid_102_to_112_v1;
wire                ready_112_to_102_v0,	ready_112_to_102_v1;
wire    [`DW-1:0]   data_112_to_122_v0,	data_112_to_122_v1;
wire                valid_112_to_122_v0,	valid_112_to_122_v1;
wire                ready_122_to_112_v0,	ready_122_to_112_v1;
wire    [`DW-1:0]   data_122_to_132_v0,	data_122_to_132_v1;
wire                valid_122_to_132_v0,	valid_122_to_132_v1;
wire                ready_132_to_122_v0,	ready_132_to_122_v1;
wire    [`DW-1:0]   data_132_to_142_v0,	data_132_to_142_v1;
wire                valid_132_to_142_v0,	valid_132_to_142_v1;
wire                ready_142_to_132_v0,	ready_142_to_132_v1;
wire    [`DW-1:0]   data_142_to_152_v0,	data_142_to_152_v1;
wire                valid_142_to_152_v0,	valid_142_to_152_v1;
wire                ready_152_to_142_v0,	ready_152_to_142_v1;
wire    [`DW-1:0]   data_152_to_162_v0,	data_152_to_162_v1;
wire                valid_152_to_162_v0,	valid_152_to_162_v1;
wire                ready_162_to_152_v0,	ready_162_to_152_v1;
wire    [`DW-1:0]   data_162_to_172_v0,	data_162_to_172_v1;
wire                valid_162_to_172_v0,	valid_162_to_172_v1;
wire                ready_172_to_162_v0,	ready_172_to_162_v1;
wire    [`DW-1:0]   data_172_to_182_v0,	data_172_to_182_v1;
wire                valid_172_to_182_v0,	valid_172_to_182_v1;
wire                ready_182_to_172_v0,	ready_182_to_172_v1;
wire    [`DW-1:0]   data_182_to_192_v0,	data_182_to_192_v1;
wire                valid_182_to_192_v0,	valid_182_to_192_v1;
wire                ready_192_to_182_v0,	ready_192_to_182_v1;
wire    [`DW-1:0]   data_192_to_202_v0,	data_192_to_202_v1;
wire                valid_192_to_202_v0,	valid_192_to_202_v1;
wire                ready_202_to_192_v0,	ready_202_to_192_v1;
wire    [`DW-1:0]   data_202_to_212_v0,	data_202_to_212_v1;
wire                valid_202_to_212_v0,	valid_202_to_212_v1;
wire                ready_212_to_202_v0,	ready_212_to_202_v1;
wire    [`DW-1:0]   data_212_to_222_v0,	data_212_to_222_v1;
wire                valid_212_to_222_v0,	valid_212_to_222_v1;
wire                ready_222_to_212_v0,	ready_222_to_212_v1;
wire    [`DW-1:0]   data_222_to_232_v0,	data_222_to_232_v1;
wire                valid_222_to_232_v0,	valid_222_to_232_v1;
wire                ready_232_to_222_v0,	ready_232_to_222_v1;
wire    [`DW-1:0]   data_232_to_242_v0,	data_232_to_242_v1;
wire                valid_232_to_242_v0,	valid_232_to_242_v1;
wire                ready_242_to_232_v0,	ready_242_to_232_v1;
wire    [`DW-1:0]   data_3_to_13_v0,	data_3_to_13_v1;
wire                valid_3_to_13_v0,	valid_3_to_13_v1;
wire                ready_13_to_3_v0,	ready_13_to_3_v1;
wire    [`DW-1:0]   data_13_to_23_v0,	data_13_to_23_v1;
wire                valid_13_to_23_v0,	valid_13_to_23_v1;
wire                ready_23_to_13_v0,	ready_23_to_13_v1;
wire    [`DW-1:0]   data_23_to_33_v0,	data_23_to_33_v1;
wire                valid_23_to_33_v0,	valid_23_to_33_v1;
wire                ready_33_to_23_v0,	ready_33_to_23_v1;
wire    [`DW-1:0]   data_33_to_43_v0,	data_33_to_43_v1;
wire                valid_33_to_43_v0,	valid_33_to_43_v1;
wire                ready_43_to_33_v0,	ready_43_to_33_v1;
wire    [`DW-1:0]   data_43_to_53_v0,	data_43_to_53_v1;
wire                valid_43_to_53_v0,	valid_43_to_53_v1;
wire                ready_53_to_43_v0,	ready_53_to_43_v1;
wire    [`DW-1:0]   data_53_to_63_v0,	data_53_to_63_v1;
wire                valid_53_to_63_v0,	valid_53_to_63_v1;
wire                ready_63_to_53_v0,	ready_63_to_53_v1;
wire    [`DW-1:0]   data_63_to_73_v0,	data_63_to_73_v1;
wire                valid_63_to_73_v0,	valid_63_to_73_v1;
wire                ready_73_to_63_v0,	ready_73_to_63_v1;
wire    [`DW-1:0]   data_73_to_83_v0,	data_73_to_83_v1;
wire                valid_73_to_83_v0,	valid_73_to_83_v1;
wire                ready_83_to_73_v0,	ready_83_to_73_v1;
wire    [`DW-1:0]   data_83_to_93_v0,	data_83_to_93_v1;
wire                valid_83_to_93_v0,	valid_83_to_93_v1;
wire                ready_93_to_83_v0,	ready_93_to_83_v1;
wire    [`DW-1:0]   data_93_to_103_v0,	data_93_to_103_v1;
wire                valid_93_to_103_v0,	valid_93_to_103_v1;
wire                ready_103_to_93_v0,	ready_103_to_93_v1;
wire    [`DW-1:0]   data_103_to_113_v0,	data_103_to_113_v1;
wire                valid_103_to_113_v0,	valid_103_to_113_v1;
wire                ready_113_to_103_v0,	ready_113_to_103_v1;
wire    [`DW-1:0]   data_113_to_123_v0,	data_113_to_123_v1;
wire                valid_113_to_123_v0,	valid_113_to_123_v1;
wire                ready_123_to_113_v0,	ready_123_to_113_v1;
wire    [`DW-1:0]   data_123_to_133_v0,	data_123_to_133_v1;
wire                valid_123_to_133_v0,	valid_123_to_133_v1;
wire                ready_133_to_123_v0,	ready_133_to_123_v1;
wire    [`DW-1:0]   data_133_to_143_v0,	data_133_to_143_v1;
wire                valid_133_to_143_v0,	valid_133_to_143_v1;
wire                ready_143_to_133_v0,	ready_143_to_133_v1;
wire    [`DW-1:0]   data_143_to_153_v0,	data_143_to_153_v1;
wire                valid_143_to_153_v0,	valid_143_to_153_v1;
wire                ready_153_to_143_v0,	ready_153_to_143_v1;
wire    [`DW-1:0]   data_153_to_163_v0,	data_153_to_163_v1;
wire                valid_153_to_163_v0,	valid_153_to_163_v1;
wire                ready_163_to_153_v0,	ready_163_to_153_v1;
wire    [`DW-1:0]   data_163_to_173_v0,	data_163_to_173_v1;
wire                valid_163_to_173_v0,	valid_163_to_173_v1;
wire                ready_173_to_163_v0,	ready_173_to_163_v1;
wire    [`DW-1:0]   data_173_to_183_v0,	data_173_to_183_v1;
wire                valid_173_to_183_v0,	valid_173_to_183_v1;
wire                ready_183_to_173_v0,	ready_183_to_173_v1;
wire    [`DW-1:0]   data_183_to_193_v0,	data_183_to_193_v1;
wire                valid_183_to_193_v0,	valid_183_to_193_v1;
wire                ready_193_to_183_v0,	ready_193_to_183_v1;
wire    [`DW-1:0]   data_193_to_203_v0,	data_193_to_203_v1;
wire                valid_193_to_203_v0,	valid_193_to_203_v1;
wire                ready_203_to_193_v0,	ready_203_to_193_v1;
wire    [`DW-1:0]   data_203_to_213_v0,	data_203_to_213_v1;
wire                valid_203_to_213_v0,	valid_203_to_213_v1;
wire                ready_213_to_203_v0,	ready_213_to_203_v1;
wire    [`DW-1:0]   data_213_to_223_v0,	data_213_to_223_v1;
wire                valid_213_to_223_v0,	valid_213_to_223_v1;
wire                ready_223_to_213_v0,	ready_223_to_213_v1;
wire    [`DW-1:0]   data_223_to_233_v0,	data_223_to_233_v1;
wire                valid_223_to_233_v0,	valid_223_to_233_v1;
wire                ready_233_to_223_v0,	ready_233_to_223_v1;
wire    [`DW-1:0]   data_233_to_243_v0,	data_233_to_243_v1;
wire                valid_233_to_243_v0,	valid_233_to_243_v1;
wire                ready_243_to_233_v0,	ready_243_to_233_v1;
wire    [`DW-1:0]   data_4_to_14_v0,	data_4_to_14_v1;
wire                valid_4_to_14_v0,	valid_4_to_14_v1;
wire                ready_14_to_4_v0,	ready_14_to_4_v1;
wire    [`DW-1:0]   data_14_to_24_v0,	data_14_to_24_v1;
wire                valid_14_to_24_v0,	valid_14_to_24_v1;
wire                ready_24_to_14_v0,	ready_24_to_14_v1;
wire    [`DW-1:0]   data_24_to_34_v0,	data_24_to_34_v1;
wire                valid_24_to_34_v0,	valid_24_to_34_v1;
wire                ready_34_to_24_v0,	ready_34_to_24_v1;
wire    [`DW-1:0]   data_34_to_44_v0,	data_34_to_44_v1;
wire                valid_34_to_44_v0,	valid_34_to_44_v1;
wire                ready_44_to_34_v0,	ready_44_to_34_v1;
wire    [`DW-1:0]   data_44_to_54_v0,	data_44_to_54_v1;
wire                valid_44_to_54_v0,	valid_44_to_54_v1;
wire                ready_54_to_44_v0,	ready_54_to_44_v1;
wire    [`DW-1:0]   data_54_to_64_v0,	data_54_to_64_v1;
wire                valid_54_to_64_v0,	valid_54_to_64_v1;
wire                ready_64_to_54_v0,	ready_64_to_54_v1;
wire    [`DW-1:0]   data_64_to_74_v0,	data_64_to_74_v1;
wire                valid_64_to_74_v0,	valid_64_to_74_v1;
wire                ready_74_to_64_v0,	ready_74_to_64_v1;
wire    [`DW-1:0]   data_74_to_84_v0,	data_74_to_84_v1;
wire                valid_74_to_84_v0,	valid_74_to_84_v1;
wire                ready_84_to_74_v0,	ready_84_to_74_v1;
wire    [`DW-1:0]   data_84_to_94_v0,	data_84_to_94_v1;
wire                valid_84_to_94_v0,	valid_84_to_94_v1;
wire                ready_94_to_84_v0,	ready_94_to_84_v1;
wire    [`DW-1:0]   data_94_to_104_v0,	data_94_to_104_v1;
wire                valid_94_to_104_v0,	valid_94_to_104_v1;
wire                ready_104_to_94_v0,	ready_104_to_94_v1;
wire    [`DW-1:0]   data_104_to_114_v0,	data_104_to_114_v1;
wire                valid_104_to_114_v0,	valid_104_to_114_v1;
wire                ready_114_to_104_v0,	ready_114_to_104_v1;
wire    [`DW-1:0]   data_114_to_124_v0,	data_114_to_124_v1;
wire                valid_114_to_124_v0,	valid_114_to_124_v1;
wire                ready_124_to_114_v0,	ready_124_to_114_v1;
wire    [`DW-1:0]   data_124_to_134_v0,	data_124_to_134_v1;
wire                valid_124_to_134_v0,	valid_124_to_134_v1;
wire                ready_134_to_124_v0,	ready_134_to_124_v1;
wire    [`DW-1:0]   data_134_to_144_v0,	data_134_to_144_v1;
wire                valid_134_to_144_v0,	valid_134_to_144_v1;
wire                ready_144_to_134_v0,	ready_144_to_134_v1;
wire    [`DW-1:0]   data_144_to_154_v0,	data_144_to_154_v1;
wire                valid_144_to_154_v0,	valid_144_to_154_v1;
wire                ready_154_to_144_v0,	ready_154_to_144_v1;
wire    [`DW-1:0]   data_154_to_164_v0,	data_154_to_164_v1;
wire                valid_154_to_164_v0,	valid_154_to_164_v1;
wire                ready_164_to_154_v0,	ready_164_to_154_v1;
wire    [`DW-1:0]   data_164_to_174_v0,	data_164_to_174_v1;
wire                valid_164_to_174_v0,	valid_164_to_174_v1;
wire                ready_174_to_164_v0,	ready_174_to_164_v1;
wire    [`DW-1:0]   data_174_to_184_v0,	data_174_to_184_v1;
wire                valid_174_to_184_v0,	valid_174_to_184_v1;
wire                ready_184_to_174_v0,	ready_184_to_174_v1;
wire    [`DW-1:0]   data_184_to_194_v0,	data_184_to_194_v1;
wire                valid_184_to_194_v0,	valid_184_to_194_v1;
wire                ready_194_to_184_v0,	ready_194_to_184_v1;
wire    [`DW-1:0]   data_194_to_204_v0,	data_194_to_204_v1;
wire                valid_194_to_204_v0,	valid_194_to_204_v1;
wire                ready_204_to_194_v0,	ready_204_to_194_v1;
wire    [`DW-1:0]   data_204_to_214_v0,	data_204_to_214_v1;
wire                valid_204_to_214_v0,	valid_204_to_214_v1;
wire                ready_214_to_204_v0,	ready_214_to_204_v1;
wire    [`DW-1:0]   data_214_to_224_v0,	data_214_to_224_v1;
wire                valid_214_to_224_v0,	valid_214_to_224_v1;
wire                ready_224_to_214_v0,	ready_224_to_214_v1;
wire    [`DW-1:0]   data_224_to_234_v0,	data_224_to_234_v1;
wire                valid_224_to_234_v0,	valid_224_to_234_v1;
wire                ready_234_to_224_v0,	ready_234_to_224_v1;
wire    [`DW-1:0]   data_234_to_244_v0,	data_234_to_244_v1;
wire                valid_234_to_244_v0,	valid_234_to_244_v1;
wire                ready_244_to_234_v0,	ready_244_to_234_v1;
wire    [`DW-1:0]   data_5_to_15_v0,	data_5_to_15_v1;
wire                valid_5_to_15_v0,	valid_5_to_15_v1;
wire                ready_15_to_5_v0,	ready_15_to_5_v1;
wire    [`DW-1:0]   data_15_to_25_v0,	data_15_to_25_v1;
wire                valid_15_to_25_v0,	valid_15_to_25_v1;
wire                ready_25_to_15_v0,	ready_25_to_15_v1;
wire    [`DW-1:0]   data_25_to_35_v0,	data_25_to_35_v1;
wire                valid_25_to_35_v0,	valid_25_to_35_v1;
wire                ready_35_to_25_v0,	ready_35_to_25_v1;
wire    [`DW-1:0]   data_35_to_45_v0,	data_35_to_45_v1;
wire                valid_35_to_45_v0,	valid_35_to_45_v1;
wire                ready_45_to_35_v0,	ready_45_to_35_v1;
wire    [`DW-1:0]   data_45_to_55_v0,	data_45_to_55_v1;
wire                valid_45_to_55_v0,	valid_45_to_55_v1;
wire                ready_55_to_45_v0,	ready_55_to_45_v1;
wire    [`DW-1:0]   data_55_to_65_v0,	data_55_to_65_v1;
wire                valid_55_to_65_v0,	valid_55_to_65_v1;
wire                ready_65_to_55_v0,	ready_65_to_55_v1;
wire    [`DW-1:0]   data_65_to_75_v0,	data_65_to_75_v1;
wire                valid_65_to_75_v0,	valid_65_to_75_v1;
wire                ready_75_to_65_v0,	ready_75_to_65_v1;
wire    [`DW-1:0]   data_75_to_85_v0,	data_75_to_85_v1;
wire                valid_75_to_85_v0,	valid_75_to_85_v1;
wire                ready_85_to_75_v0,	ready_85_to_75_v1;
wire    [`DW-1:0]   data_85_to_95_v0,	data_85_to_95_v1;
wire                valid_85_to_95_v0,	valid_85_to_95_v1;
wire                ready_95_to_85_v0,	ready_95_to_85_v1;
wire    [`DW-1:0]   data_95_to_105_v0,	data_95_to_105_v1;
wire                valid_95_to_105_v0,	valid_95_to_105_v1;
wire                ready_105_to_95_v0,	ready_105_to_95_v1;
wire    [`DW-1:0]   data_105_to_115_v0,	data_105_to_115_v1;
wire                valid_105_to_115_v0,	valid_105_to_115_v1;
wire                ready_115_to_105_v0,	ready_115_to_105_v1;
wire    [`DW-1:0]   data_115_to_125_v0,	data_115_to_125_v1;
wire                valid_115_to_125_v0,	valid_115_to_125_v1;
wire                ready_125_to_115_v0,	ready_125_to_115_v1;
wire    [`DW-1:0]   data_125_to_135_v0,	data_125_to_135_v1;
wire                valid_125_to_135_v0,	valid_125_to_135_v1;
wire                ready_135_to_125_v0,	ready_135_to_125_v1;
wire    [`DW-1:0]   data_135_to_145_v0,	data_135_to_145_v1;
wire                valid_135_to_145_v0,	valid_135_to_145_v1;
wire                ready_145_to_135_v0,	ready_145_to_135_v1;
wire    [`DW-1:0]   data_145_to_155_v0,	data_145_to_155_v1;
wire                valid_145_to_155_v0,	valid_145_to_155_v1;
wire                ready_155_to_145_v0,	ready_155_to_145_v1;
wire    [`DW-1:0]   data_155_to_165_v0,	data_155_to_165_v1;
wire                valid_155_to_165_v0,	valid_155_to_165_v1;
wire                ready_165_to_155_v0,	ready_165_to_155_v1;
wire    [`DW-1:0]   data_165_to_175_v0,	data_165_to_175_v1;
wire                valid_165_to_175_v0,	valid_165_to_175_v1;
wire                ready_175_to_165_v0,	ready_175_to_165_v1;
wire    [`DW-1:0]   data_175_to_185_v0,	data_175_to_185_v1;
wire                valid_175_to_185_v0,	valid_175_to_185_v1;
wire                ready_185_to_175_v0,	ready_185_to_175_v1;
wire    [`DW-1:0]   data_185_to_195_v0,	data_185_to_195_v1;
wire                valid_185_to_195_v0,	valid_185_to_195_v1;
wire                ready_195_to_185_v0,	ready_195_to_185_v1;
wire    [`DW-1:0]   data_195_to_205_v0,	data_195_to_205_v1;
wire                valid_195_to_205_v0,	valid_195_to_205_v1;
wire                ready_205_to_195_v0,	ready_205_to_195_v1;
wire    [`DW-1:0]   data_205_to_215_v0,	data_205_to_215_v1;
wire                valid_205_to_215_v0,	valid_205_to_215_v1;
wire                ready_215_to_205_v0,	ready_215_to_205_v1;
wire    [`DW-1:0]   data_215_to_225_v0,	data_215_to_225_v1;
wire                valid_215_to_225_v0,	valid_215_to_225_v1;
wire                ready_225_to_215_v0,	ready_225_to_215_v1;
wire    [`DW-1:0]   data_225_to_235_v0,	data_225_to_235_v1;
wire                valid_225_to_235_v0,	valid_225_to_235_v1;
wire                ready_235_to_225_v0,	ready_235_to_225_v1;
wire    [`DW-1:0]   data_235_to_245_v0,	data_235_to_245_v1;
wire                valid_235_to_245_v0,	valid_235_to_245_v1;
wire                ready_245_to_235_v0,	ready_245_to_235_v1;
wire    [`DW-1:0]   data_6_to_16_v0,	data_6_to_16_v1;
wire                valid_6_to_16_v0,	valid_6_to_16_v1;
wire                ready_16_to_6_v0,	ready_16_to_6_v1;
wire    [`DW-1:0]   data_16_to_26_v0,	data_16_to_26_v1;
wire                valid_16_to_26_v0,	valid_16_to_26_v1;
wire                ready_26_to_16_v0,	ready_26_to_16_v1;
wire    [`DW-1:0]   data_26_to_36_v0,	data_26_to_36_v1;
wire                valid_26_to_36_v0,	valid_26_to_36_v1;
wire                ready_36_to_26_v0,	ready_36_to_26_v1;
wire    [`DW-1:0]   data_36_to_46_v0,	data_36_to_46_v1;
wire                valid_36_to_46_v0,	valid_36_to_46_v1;
wire                ready_46_to_36_v0,	ready_46_to_36_v1;
wire    [`DW-1:0]   data_46_to_56_v0,	data_46_to_56_v1;
wire                valid_46_to_56_v0,	valid_46_to_56_v1;
wire                ready_56_to_46_v0,	ready_56_to_46_v1;
wire    [`DW-1:0]   data_56_to_66_v0,	data_56_to_66_v1;
wire                valid_56_to_66_v0,	valid_56_to_66_v1;
wire                ready_66_to_56_v0,	ready_66_to_56_v1;
wire    [`DW-1:0]   data_66_to_76_v0,	data_66_to_76_v1;
wire                valid_66_to_76_v0,	valid_66_to_76_v1;
wire                ready_76_to_66_v0,	ready_76_to_66_v1;
wire    [`DW-1:0]   data_76_to_86_v0,	data_76_to_86_v1;
wire                valid_76_to_86_v0,	valid_76_to_86_v1;
wire                ready_86_to_76_v0,	ready_86_to_76_v1;
wire    [`DW-1:0]   data_86_to_96_v0,	data_86_to_96_v1;
wire                valid_86_to_96_v0,	valid_86_to_96_v1;
wire                ready_96_to_86_v0,	ready_96_to_86_v1;
wire    [`DW-1:0]   data_96_to_106_v0,	data_96_to_106_v1;
wire                valid_96_to_106_v0,	valid_96_to_106_v1;
wire                ready_106_to_96_v0,	ready_106_to_96_v1;
wire    [`DW-1:0]   data_106_to_116_v0,	data_106_to_116_v1;
wire                valid_106_to_116_v0,	valid_106_to_116_v1;
wire                ready_116_to_106_v0,	ready_116_to_106_v1;
wire    [`DW-1:0]   data_116_to_126_v0,	data_116_to_126_v1;
wire                valid_116_to_126_v0,	valid_116_to_126_v1;
wire                ready_126_to_116_v0,	ready_126_to_116_v1;
wire    [`DW-1:0]   data_126_to_136_v0,	data_126_to_136_v1;
wire                valid_126_to_136_v0,	valid_126_to_136_v1;
wire                ready_136_to_126_v0,	ready_136_to_126_v1;
wire    [`DW-1:0]   data_136_to_146_v0,	data_136_to_146_v1;
wire                valid_136_to_146_v0,	valid_136_to_146_v1;
wire                ready_146_to_136_v0,	ready_146_to_136_v1;
wire    [`DW-1:0]   data_146_to_156_v0,	data_146_to_156_v1;
wire                valid_146_to_156_v0,	valid_146_to_156_v1;
wire                ready_156_to_146_v0,	ready_156_to_146_v1;
wire    [`DW-1:0]   data_156_to_166_v0,	data_156_to_166_v1;
wire                valid_156_to_166_v0,	valid_156_to_166_v1;
wire                ready_166_to_156_v0,	ready_166_to_156_v1;
wire    [`DW-1:0]   data_166_to_176_v0,	data_166_to_176_v1;
wire                valid_166_to_176_v0,	valid_166_to_176_v1;
wire                ready_176_to_166_v0,	ready_176_to_166_v1;
wire    [`DW-1:0]   data_176_to_186_v0,	data_176_to_186_v1;
wire                valid_176_to_186_v0,	valid_176_to_186_v1;
wire                ready_186_to_176_v0,	ready_186_to_176_v1;
wire    [`DW-1:0]   data_186_to_196_v0,	data_186_to_196_v1;
wire                valid_186_to_196_v0,	valid_186_to_196_v1;
wire                ready_196_to_186_v0,	ready_196_to_186_v1;
wire    [`DW-1:0]   data_196_to_206_v0,	data_196_to_206_v1;
wire                valid_196_to_206_v0,	valid_196_to_206_v1;
wire                ready_206_to_196_v0,	ready_206_to_196_v1;
wire    [`DW-1:0]   data_206_to_216_v0,	data_206_to_216_v1;
wire                valid_206_to_216_v0,	valid_206_to_216_v1;
wire                ready_216_to_206_v0,	ready_216_to_206_v1;
wire    [`DW-1:0]   data_216_to_226_v0,	data_216_to_226_v1;
wire                valid_216_to_226_v0,	valid_216_to_226_v1;
wire                ready_226_to_216_v0,	ready_226_to_216_v1;
wire    [`DW-1:0]   data_226_to_236_v0,	data_226_to_236_v1;
wire                valid_226_to_236_v0,	valid_226_to_236_v1;
wire                ready_236_to_226_v0,	ready_236_to_226_v1;
wire    [`DW-1:0]   data_236_to_246_v0,	data_236_to_246_v1;
wire                valid_236_to_246_v0,	valid_236_to_246_v1;
wire                ready_246_to_236_v0,	ready_246_to_236_v1;
wire    [`DW-1:0]   data_7_to_17_v0,	data_7_to_17_v1;
wire                valid_7_to_17_v0,	valid_7_to_17_v1;
wire                ready_17_to_7_v0,	ready_17_to_7_v1;
wire    [`DW-1:0]   data_17_to_27_v0,	data_17_to_27_v1;
wire                valid_17_to_27_v0,	valid_17_to_27_v1;
wire                ready_27_to_17_v0,	ready_27_to_17_v1;
wire    [`DW-1:0]   data_27_to_37_v0,	data_27_to_37_v1;
wire                valid_27_to_37_v0,	valid_27_to_37_v1;
wire                ready_37_to_27_v0,	ready_37_to_27_v1;
wire    [`DW-1:0]   data_37_to_47_v0,	data_37_to_47_v1;
wire                valid_37_to_47_v0,	valid_37_to_47_v1;
wire                ready_47_to_37_v0,	ready_47_to_37_v1;
wire    [`DW-1:0]   data_47_to_57_v0,	data_47_to_57_v1;
wire                valid_47_to_57_v0,	valid_47_to_57_v1;
wire                ready_57_to_47_v0,	ready_57_to_47_v1;
wire    [`DW-1:0]   data_57_to_67_v0,	data_57_to_67_v1;
wire                valid_57_to_67_v0,	valid_57_to_67_v1;
wire                ready_67_to_57_v0,	ready_67_to_57_v1;
wire    [`DW-1:0]   data_67_to_77_v0,	data_67_to_77_v1;
wire                valid_67_to_77_v0,	valid_67_to_77_v1;
wire                ready_77_to_67_v0,	ready_77_to_67_v1;
wire    [`DW-1:0]   data_77_to_87_v0,	data_77_to_87_v1;
wire                valid_77_to_87_v0,	valid_77_to_87_v1;
wire                ready_87_to_77_v0,	ready_87_to_77_v1;
wire    [`DW-1:0]   data_87_to_97_v0,	data_87_to_97_v1;
wire                valid_87_to_97_v0,	valid_87_to_97_v1;
wire                ready_97_to_87_v0,	ready_97_to_87_v1;
wire    [`DW-1:0]   data_97_to_107_v0,	data_97_to_107_v1;
wire                valid_97_to_107_v0,	valid_97_to_107_v1;
wire                ready_107_to_97_v0,	ready_107_to_97_v1;
wire    [`DW-1:0]   data_107_to_117_v0,	data_107_to_117_v1;
wire                valid_107_to_117_v0,	valid_107_to_117_v1;
wire                ready_117_to_107_v0,	ready_117_to_107_v1;
wire    [`DW-1:0]   data_117_to_127_v0,	data_117_to_127_v1;
wire                valid_117_to_127_v0,	valid_117_to_127_v1;
wire                ready_127_to_117_v0,	ready_127_to_117_v1;
wire    [`DW-1:0]   data_127_to_137_v0,	data_127_to_137_v1;
wire                valid_127_to_137_v0,	valid_127_to_137_v1;
wire                ready_137_to_127_v0,	ready_137_to_127_v1;
wire    [`DW-1:0]   data_137_to_147_v0,	data_137_to_147_v1;
wire                valid_137_to_147_v0,	valid_137_to_147_v1;
wire                ready_147_to_137_v0,	ready_147_to_137_v1;
wire    [`DW-1:0]   data_147_to_157_v0,	data_147_to_157_v1;
wire                valid_147_to_157_v0,	valid_147_to_157_v1;
wire                ready_157_to_147_v0,	ready_157_to_147_v1;
wire    [`DW-1:0]   data_157_to_167_v0,	data_157_to_167_v1;
wire                valid_157_to_167_v0,	valid_157_to_167_v1;
wire                ready_167_to_157_v0,	ready_167_to_157_v1;
wire    [`DW-1:0]   data_167_to_177_v0,	data_167_to_177_v1;
wire                valid_167_to_177_v0,	valid_167_to_177_v1;
wire                ready_177_to_167_v0,	ready_177_to_167_v1;
wire    [`DW-1:0]   data_177_to_187_v0,	data_177_to_187_v1;
wire                valid_177_to_187_v0,	valid_177_to_187_v1;
wire                ready_187_to_177_v0,	ready_187_to_177_v1;
wire    [`DW-1:0]   data_187_to_197_v0,	data_187_to_197_v1;
wire                valid_187_to_197_v0,	valid_187_to_197_v1;
wire                ready_197_to_187_v0,	ready_197_to_187_v1;
wire    [`DW-1:0]   data_197_to_207_v0,	data_197_to_207_v1;
wire                valid_197_to_207_v0,	valid_197_to_207_v1;
wire                ready_207_to_197_v0,	ready_207_to_197_v1;
wire    [`DW-1:0]   data_207_to_217_v0,	data_207_to_217_v1;
wire                valid_207_to_217_v0,	valid_207_to_217_v1;
wire                ready_217_to_207_v0,	ready_217_to_207_v1;
wire    [`DW-1:0]   data_217_to_227_v0,	data_217_to_227_v1;
wire                valid_217_to_227_v0,	valid_217_to_227_v1;
wire                ready_227_to_217_v0,	ready_227_to_217_v1;
wire    [`DW-1:0]   data_227_to_237_v0,	data_227_to_237_v1;
wire                valid_227_to_237_v0,	valid_227_to_237_v1;
wire                ready_237_to_227_v0,	ready_237_to_227_v1;
wire    [`DW-1:0]   data_237_to_247_v0,	data_237_to_247_v1;
wire                valid_237_to_247_v0,	valid_237_to_247_v1;
wire                ready_247_to_237_v0,	ready_247_to_237_v1;
wire    [`DW-1:0]   data_8_to_18_v0,	data_8_to_18_v1;
wire                valid_8_to_18_v0,	valid_8_to_18_v1;
wire                ready_18_to_8_v0,	ready_18_to_8_v1;
wire    [`DW-1:0]   data_18_to_28_v0,	data_18_to_28_v1;
wire                valid_18_to_28_v0,	valid_18_to_28_v1;
wire                ready_28_to_18_v0,	ready_28_to_18_v1;
wire    [`DW-1:0]   data_28_to_38_v0,	data_28_to_38_v1;
wire                valid_28_to_38_v0,	valid_28_to_38_v1;
wire                ready_38_to_28_v0,	ready_38_to_28_v1;
wire    [`DW-1:0]   data_38_to_48_v0,	data_38_to_48_v1;
wire                valid_38_to_48_v0,	valid_38_to_48_v1;
wire                ready_48_to_38_v0,	ready_48_to_38_v1;
wire    [`DW-1:0]   data_48_to_58_v0,	data_48_to_58_v1;
wire                valid_48_to_58_v0,	valid_48_to_58_v1;
wire                ready_58_to_48_v0,	ready_58_to_48_v1;
wire    [`DW-1:0]   data_58_to_68_v0,	data_58_to_68_v1;
wire                valid_58_to_68_v0,	valid_58_to_68_v1;
wire                ready_68_to_58_v0,	ready_68_to_58_v1;
wire    [`DW-1:0]   data_68_to_78_v0,	data_68_to_78_v1;
wire                valid_68_to_78_v0,	valid_68_to_78_v1;
wire                ready_78_to_68_v0,	ready_78_to_68_v1;
wire    [`DW-1:0]   data_78_to_88_v0,	data_78_to_88_v1;
wire                valid_78_to_88_v0,	valid_78_to_88_v1;
wire                ready_88_to_78_v0,	ready_88_to_78_v1;
wire    [`DW-1:0]   data_88_to_98_v0,	data_88_to_98_v1;
wire                valid_88_to_98_v0,	valid_88_to_98_v1;
wire                ready_98_to_88_v0,	ready_98_to_88_v1;
wire    [`DW-1:0]   data_98_to_108_v0,	data_98_to_108_v1;
wire                valid_98_to_108_v0,	valid_98_to_108_v1;
wire                ready_108_to_98_v0,	ready_108_to_98_v1;
wire    [`DW-1:0]   data_108_to_118_v0,	data_108_to_118_v1;
wire                valid_108_to_118_v0,	valid_108_to_118_v1;
wire                ready_118_to_108_v0,	ready_118_to_108_v1;
wire    [`DW-1:0]   data_118_to_128_v0,	data_118_to_128_v1;
wire                valid_118_to_128_v0,	valid_118_to_128_v1;
wire                ready_128_to_118_v0,	ready_128_to_118_v1;
wire    [`DW-1:0]   data_128_to_138_v0,	data_128_to_138_v1;
wire                valid_128_to_138_v0,	valid_128_to_138_v1;
wire                ready_138_to_128_v0,	ready_138_to_128_v1;
wire    [`DW-1:0]   data_138_to_148_v0,	data_138_to_148_v1;
wire                valid_138_to_148_v0,	valid_138_to_148_v1;
wire                ready_148_to_138_v0,	ready_148_to_138_v1;
wire    [`DW-1:0]   data_148_to_158_v0,	data_148_to_158_v1;
wire                valid_148_to_158_v0,	valid_148_to_158_v1;
wire                ready_158_to_148_v0,	ready_158_to_148_v1;
wire    [`DW-1:0]   data_158_to_168_v0,	data_158_to_168_v1;
wire                valid_158_to_168_v0,	valid_158_to_168_v1;
wire                ready_168_to_158_v0,	ready_168_to_158_v1;
wire    [`DW-1:0]   data_168_to_178_v0,	data_168_to_178_v1;
wire                valid_168_to_178_v0,	valid_168_to_178_v1;
wire                ready_178_to_168_v0,	ready_178_to_168_v1;
wire    [`DW-1:0]   data_178_to_188_v0,	data_178_to_188_v1;
wire                valid_178_to_188_v0,	valid_178_to_188_v1;
wire                ready_188_to_178_v0,	ready_188_to_178_v1;
wire    [`DW-1:0]   data_188_to_198_v0,	data_188_to_198_v1;
wire                valid_188_to_198_v0,	valid_188_to_198_v1;
wire                ready_198_to_188_v0,	ready_198_to_188_v1;
wire    [`DW-1:0]   data_198_to_208_v0,	data_198_to_208_v1;
wire                valid_198_to_208_v0,	valid_198_to_208_v1;
wire                ready_208_to_198_v0,	ready_208_to_198_v1;
wire    [`DW-1:0]   data_208_to_218_v0,	data_208_to_218_v1;
wire                valid_208_to_218_v0,	valid_208_to_218_v1;
wire                ready_218_to_208_v0,	ready_218_to_208_v1;
wire    [`DW-1:0]   data_218_to_228_v0,	data_218_to_228_v1;
wire                valid_218_to_228_v0,	valid_218_to_228_v1;
wire                ready_228_to_218_v0,	ready_228_to_218_v1;
wire    [`DW-1:0]   data_228_to_238_v0,	data_228_to_238_v1;
wire                valid_228_to_238_v0,	valid_228_to_238_v1;
wire                ready_238_to_228_v0,	ready_238_to_228_v1;
wire    [`DW-1:0]   data_238_to_248_v0,	data_238_to_248_v1;
wire                valid_238_to_248_v0,	valid_238_to_248_v1;
wire                ready_248_to_238_v0,	ready_248_to_238_v1;
wire    [`DW-1:0]   data_9_to_19_v0,	data_9_to_19_v1;
wire                valid_9_to_19_v0,	valid_9_to_19_v1;
wire                ready_19_to_9_v0,	ready_19_to_9_v1;
wire    [`DW-1:0]   data_19_to_29_v0,	data_19_to_29_v1;
wire                valid_19_to_29_v0,	valid_19_to_29_v1;
wire                ready_29_to_19_v0,	ready_29_to_19_v1;
wire    [`DW-1:0]   data_29_to_39_v0,	data_29_to_39_v1;
wire                valid_29_to_39_v0,	valid_29_to_39_v1;
wire                ready_39_to_29_v0,	ready_39_to_29_v1;
wire    [`DW-1:0]   data_39_to_49_v0,	data_39_to_49_v1;
wire                valid_39_to_49_v0,	valid_39_to_49_v1;
wire                ready_49_to_39_v0,	ready_49_to_39_v1;
wire    [`DW-1:0]   data_49_to_59_v0,	data_49_to_59_v1;
wire                valid_49_to_59_v0,	valid_49_to_59_v1;
wire                ready_59_to_49_v0,	ready_59_to_49_v1;
wire    [`DW-1:0]   data_59_to_69_v0,	data_59_to_69_v1;
wire                valid_59_to_69_v0,	valid_59_to_69_v1;
wire                ready_69_to_59_v0,	ready_69_to_59_v1;
wire    [`DW-1:0]   data_69_to_79_v0,	data_69_to_79_v1;
wire                valid_69_to_79_v0,	valid_69_to_79_v1;
wire                ready_79_to_69_v0,	ready_79_to_69_v1;
wire    [`DW-1:0]   data_79_to_89_v0,	data_79_to_89_v1;
wire                valid_79_to_89_v0,	valid_79_to_89_v1;
wire                ready_89_to_79_v0,	ready_89_to_79_v1;
wire    [`DW-1:0]   data_89_to_99_v0,	data_89_to_99_v1;
wire                valid_89_to_99_v0,	valid_89_to_99_v1;
wire                ready_99_to_89_v0,	ready_99_to_89_v1;
wire    [`DW-1:0]   data_99_to_109_v0,	data_99_to_109_v1;
wire                valid_99_to_109_v0,	valid_99_to_109_v1;
wire                ready_109_to_99_v0,	ready_109_to_99_v1;
wire    [`DW-1:0]   data_109_to_119_v0,	data_109_to_119_v1;
wire                valid_109_to_119_v0,	valid_109_to_119_v1;
wire                ready_119_to_109_v0,	ready_119_to_109_v1;
wire    [`DW-1:0]   data_119_to_129_v0,	data_119_to_129_v1;
wire                valid_119_to_129_v0,	valid_119_to_129_v1;
wire                ready_129_to_119_v0,	ready_129_to_119_v1;
wire    [`DW-1:0]   data_129_to_139_v0,	data_129_to_139_v1;
wire                valid_129_to_139_v0,	valid_129_to_139_v1;
wire                ready_139_to_129_v0,	ready_139_to_129_v1;
wire    [`DW-1:0]   data_139_to_149_v0,	data_139_to_149_v1;
wire                valid_139_to_149_v0,	valid_139_to_149_v1;
wire                ready_149_to_139_v0,	ready_149_to_139_v1;
wire    [`DW-1:0]   data_149_to_159_v0,	data_149_to_159_v1;
wire                valid_149_to_159_v0,	valid_149_to_159_v1;
wire                ready_159_to_149_v0,	ready_159_to_149_v1;
wire    [`DW-1:0]   data_159_to_169_v0,	data_159_to_169_v1;
wire                valid_159_to_169_v0,	valid_159_to_169_v1;
wire                ready_169_to_159_v0,	ready_169_to_159_v1;
wire    [`DW-1:0]   data_169_to_179_v0,	data_169_to_179_v1;
wire                valid_169_to_179_v0,	valid_169_to_179_v1;
wire                ready_179_to_169_v0,	ready_179_to_169_v1;
wire    [`DW-1:0]   data_179_to_189_v0,	data_179_to_189_v1;
wire                valid_179_to_189_v0,	valid_179_to_189_v1;
wire                ready_189_to_179_v0,	ready_189_to_179_v1;
wire    [`DW-1:0]   data_189_to_199_v0,	data_189_to_199_v1;
wire                valid_189_to_199_v0,	valid_189_to_199_v1;
wire                ready_199_to_189_v0,	ready_199_to_189_v1;
wire    [`DW-1:0]   data_199_to_209_v0,	data_199_to_209_v1;
wire                valid_199_to_209_v0,	valid_199_to_209_v1;
wire                ready_209_to_199_v0,	ready_209_to_199_v1;
wire    [`DW-1:0]   data_209_to_219_v0,	data_209_to_219_v1;
wire                valid_209_to_219_v0,	valid_209_to_219_v1;
wire                ready_219_to_209_v0,	ready_219_to_209_v1;
wire    [`DW-1:0]   data_219_to_229_v0,	data_219_to_229_v1;
wire                valid_219_to_229_v0,	valid_219_to_229_v1;
wire                ready_229_to_219_v0,	ready_229_to_219_v1;
wire    [`DW-1:0]   data_229_to_239_v0,	data_229_to_239_v1;
wire                valid_229_to_239_v0,	valid_229_to_239_v1;
wire                ready_239_to_229_v0,	ready_239_to_229_v1;
wire    [`DW-1:0]   data_239_to_249_v0,	data_239_to_249_v1;
wire                valid_239_to_249_v0,	valid_239_to_249_v1;
wire                ready_249_to_239_v0,	ready_249_to_239_v1;

/*Router 0,0*/    
cast_router #(
    .isUBM_list            (isUBM_list_0_0),
    .isFC_list             (isFC_list_0_0),
    .FCdn_list             (FCdn_list_0_0),
    .FCpl_list             (FCpl_list_0_0),
    .rt_file_list          (cast_rt_file_list_0_0)
)router_0_0(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_i_stab),
    .west_valid_i          (valid_i_stab),
    .west_ready_o          (ready_o_stab),
    .west_data_o           (),
    .west_valid_o          (),
    .west_ready_i          (1'b0),
    .east_data_i           (data_1_to_0),
    .east_valid_i          (valid_1_to_0),
    .east_ready_o          (ready_0_to_1),
    .east_data_o           (data_0_to_1),
    .east_valid_o          (valid_0_to_1),
    .east_ready_i          (ready_1_to_0),
    .vert0_data_i          (34'b0),
    .vert0_valid_i         (1'b0),
    .vert0_ready_o         (),
    .vert0_data_o          (data_0_to_10_v0),
    .vert0_valid_o         (valid_0_to_10_v0),
    .vert0_ready_i         (ready_10_to_0_v0),
    .vert1_data_i          (34'b0),
    .vert1_valid_i         (1'b0),
    .vert1_ready_o         (),
    .vert1_data_o          (data_0_to_10_v1),
    .vert1_valid_o         (valid_0_to_10_v1),
    .vert1_ready_i         (ready_10_to_0_v1),
    .local_data_i          (data_i[0][0]),
    .local_valid_i         (valid_i[0][0]),
    .local_ready_o         (ready_o[0][0]),
    .local_data_o          (data_o[0][0]),
    .local_valid_o         (valid_o[0][0]),
    .local_ready_i         (ready_i[0][0]),
    .credit_upd            (credit_upd)
);

/*Router 0,1*/    
cast_router #(
    .isUBM_list            (isUBM_list_0_1),
    .isFC_list             (isFC_list_0_1),
    .FCdn_list             (FCdn_list_0_1),
    .FCpl_list             (FCpl_list_0_1),
    .rt_file_list          (cast_rt_file_list_0_1)
)router_0_1(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (34'b0),
    .west_valid_i          (1'b0),
    .west_ready_o          (),
    .west_data_o           (),
    .west_valid_o          (),
    .west_ready_i          (1'b0),
    .east_data_i           (data_11_to_10),
    .east_valid_i          (valid_11_to_10),
    .east_ready_o          (ready_10_to_11),
    .east_data_o           (data_10_to_11),
    .east_valid_o          (valid_10_to_11),
    .east_ready_i          (ready_11_to_10),
    .vert0_data_i          (data_0_to_10_v0),
    .vert0_valid_i         (valid_0_to_10_v0),
    .vert0_ready_o         (ready_10_to_0_v0),
    .vert0_data_o          (data_10_to_20_v0),
    .vert0_valid_o         (valid_10_to_20_v0),
    .vert0_ready_i         (ready_20_to_10_v0),
    .vert1_data_i          (data_0_to_10_v1),
    .vert1_valid_i         (valid_0_to_10_v1),
    .vert1_ready_o         (ready_10_to_0_v1),
    .vert1_data_o          (data_10_to_20_v1),
    .vert1_valid_o         (valid_10_to_20_v1),
    .vert1_ready_i         (ready_20_to_10_v1),
    .local_data_i          (data_i[0][1]),
    .local_valid_i         (valid_i[0][1]),
    .local_ready_o         (ready_o[0][1]),
    .local_data_o          (data_o[0][1]),
    .local_valid_o         (valid_o[0][1]),
    .local_ready_i         (ready_i[0][1]),
    .credit_upd            (credit_upd)
);

/*Router 0,2*/    
cast_router #(
    .isUBM_list            (isUBM_list_0_2),
    .isFC_list             (isFC_list_0_2),
    .FCdn_list             (FCdn_list_0_2),
    .FCpl_list             (FCpl_list_0_2),
    .rt_file_list          (cast_rt_file_list_0_2)
)router_0_2(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (34'b0),
    .west_valid_i          (1'b0),
    .west_ready_o          (),
    .west_data_o           (),
    .west_valid_o          (),
    .west_ready_i          (1'b0),
    .east_data_i           (data_21_to_20),
    .east_valid_i          (valid_21_to_20),
    .east_ready_o          (ready_20_to_21),
    .east_data_o           (data_20_to_21),
    .east_valid_o          (valid_20_to_21),
    .east_ready_i          (ready_21_to_20),
    .vert0_data_i          (data_10_to_20_v0),
    .vert0_valid_i         (valid_10_to_20_v0),
    .vert0_ready_o         (ready_20_to_10_v0),
    .vert0_data_o          (data_20_to_30_v0),
    .vert0_valid_o         (valid_20_to_30_v0),
    .vert0_ready_i         (ready_30_to_20_v0),
    .vert1_data_i          (data_10_to_20_v1),
    .vert1_valid_i         (valid_10_to_20_v1),
    .vert1_ready_o         (ready_20_to_10_v1),
    .vert1_data_o          (data_20_to_30_v1),
    .vert1_valid_o         (valid_20_to_30_v1),
    .vert1_ready_i         (ready_30_to_20_v1),
    .local_data_i          (data_i[0][2]),
    .local_valid_i         (valid_i[0][2]),
    .local_ready_o         (ready_o[0][2]),
    .local_data_o          (data_o[0][2]),
    .local_valid_o         (valid_o[0][2]),
    .local_ready_i         (ready_i[0][2]),
    .credit_upd            (credit_upd)
);

/*Router 0,3*/    
cast_router #(
    .isUBM_list            (isUBM_list_0_3),
    .isFC_list             (isFC_list_0_3),
    .FCdn_list             (FCdn_list_0_3),
    .FCpl_list             (FCpl_list_0_3),
    .rt_file_list          (cast_rt_file_list_0_3)
)router_0_3(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (34'b0),
    .west_valid_i          (1'b0),
    .west_ready_o          (),
    .west_data_o           (),
    .west_valid_o          (),
    .west_ready_i          (1'b0),
    .east_data_i           (data_31_to_30),
    .east_valid_i          (valid_31_to_30),
    .east_ready_o          (ready_30_to_31),
    .east_data_o           (data_30_to_31),
    .east_valid_o          (valid_30_to_31),
    .east_ready_i          (ready_31_to_30),
    .vert0_data_i          (data_20_to_30_v0),
    .vert0_valid_i         (valid_20_to_30_v0),
    .vert0_ready_o         (ready_30_to_20_v0),
    .vert0_data_o          (data_30_to_40_v0),
    .vert0_valid_o         (valid_30_to_40_v0),
    .vert0_ready_i         (ready_40_to_30_v0),
    .vert1_data_i          (data_20_to_30_v1),
    .vert1_valid_i         (valid_20_to_30_v1),
    .vert1_ready_o         (ready_30_to_20_v1),
    .vert1_data_o          (data_30_to_40_v1),
    .vert1_valid_o         (valid_30_to_40_v1),
    .vert1_ready_i         (ready_40_to_30_v1),
    .local_data_i          (data_i[0][3]),
    .local_valid_i         (valid_i[0][3]),
    .local_ready_o         (ready_o[0][3]),
    .local_data_o          (data_o[0][3]),
    .local_valid_o         (valid_o[0][3]),
    .local_ready_i         (ready_i[0][3]),
    .credit_upd            (credit_upd)
);

/*Router 0,4*/    
cast_router #(
    .isUBM_list            (isUBM_list_0_4),
    .isFC_list             (isFC_list_0_4),
    .FCdn_list             (FCdn_list_0_4),
    .FCpl_list             (FCpl_list_0_4),
    .rt_file_list          (cast_rt_file_list_0_4)
)router_0_4(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (34'b0),
    .west_valid_i          (1'b0),
    .west_ready_o          (),
    .west_data_o           (),
    .west_valid_o          (),
    .west_ready_i          (1'b0),
    .east_data_i           (data_41_to_40),
    .east_valid_i          (valid_41_to_40),
    .east_ready_o          (ready_40_to_41),
    .east_data_o           (data_40_to_41),
    .east_valid_o          (valid_40_to_41),
    .east_ready_i          (ready_41_to_40),
    .vert0_data_i          (data_30_to_40_v0),
    .vert0_valid_i         (valid_30_to_40_v0),
    .vert0_ready_o         (ready_40_to_30_v0),
    .vert0_data_o          (data_40_to_50_v0),
    .vert0_valid_o         (valid_40_to_50_v0),
    .vert0_ready_i         (ready_50_to_40_v0),
    .vert1_data_i          (data_30_to_40_v1),
    .vert1_valid_i         (valid_30_to_40_v1),
    .vert1_ready_o         (ready_40_to_30_v1),
    .vert1_data_o          (data_40_to_50_v1),
    .vert1_valid_o         (valid_40_to_50_v1),
    .vert1_ready_i         (ready_50_to_40_v1),
    .local_data_i          (data_i[0][4]),
    .local_valid_i         (valid_i[0][4]),
    .local_ready_o         (ready_o[0][4]),
    .local_data_o          (data_o[0][4]),
    .local_valid_o         (valid_o[0][4]),
    .local_ready_i         (ready_i[0][4]),
    .credit_upd            (credit_upd)
);

/*Router 0,5*/    
cast_router #(
    .isUBM_list            (isUBM_list_0_5),
    .isFC_list             (isFC_list_0_5),
    .FCdn_list             (FCdn_list_0_5),
    .FCpl_list             (FCpl_list_0_5),
    .rt_file_list          (cast_rt_file_list_0_5)
)router_0_5(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (34'b0),
    .west_valid_i          (1'b0),
    .west_ready_o          (),
    .west_data_o           (),
    .west_valid_o          (),
    .west_ready_i          (1'b0),
    .east_data_i           (data_51_to_50),
    .east_valid_i          (valid_51_to_50),
    .east_ready_o          (ready_50_to_51),
    .east_data_o           (data_50_to_51),
    .east_valid_o          (valid_50_to_51),
    .east_ready_i          (ready_51_to_50),
    .vert0_data_i          (data_40_to_50_v0),
    .vert0_valid_i         (valid_40_to_50_v0),
    .vert0_ready_o         (ready_50_to_40_v0),
    .vert0_data_o          (data_50_to_60_v0),
    .vert0_valid_o         (valid_50_to_60_v0),
    .vert0_ready_i         (ready_60_to_50_v0),
    .vert1_data_i          (data_40_to_50_v1),
    .vert1_valid_i         (valid_40_to_50_v1),
    .vert1_ready_o         (ready_50_to_40_v1),
    .vert1_data_o          (data_50_to_60_v1),
    .vert1_valid_o         (valid_50_to_60_v1),
    .vert1_ready_i         (ready_60_to_50_v1),
    .local_data_i          (data_i[0][5]),
    .local_valid_i         (valid_i[0][5]),
    .local_ready_o         (ready_o[0][5]),
    .local_data_o          (data_o[0][5]),
    .local_valid_o         (valid_o[0][5]),
    .local_ready_i         (ready_i[0][5]),
    .credit_upd            (credit_upd)
);

/*Router 0,6*/    
cast_router #(
    .isUBM_list            (isUBM_list_0_6),
    .isFC_list             (isFC_list_0_6),
    .FCdn_list             (FCdn_list_0_6),
    .FCpl_list             (FCpl_list_0_6),
    .rt_file_list          (cast_rt_file_list_0_6)
)router_0_6(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (34'b0),
    .west_valid_i          (1'b0),
    .west_ready_o          (),
    .west_data_o           (),
    .west_valid_o          (),
    .west_ready_i          (1'b0),
    .east_data_i           (data_61_to_60),
    .east_valid_i          (valid_61_to_60),
    .east_ready_o          (ready_60_to_61),
    .east_data_o           (data_60_to_61),
    .east_valid_o          (valid_60_to_61),
    .east_ready_i          (ready_61_to_60),
    .vert0_data_i          (data_50_to_60_v0),
    .vert0_valid_i         (valid_50_to_60_v0),
    .vert0_ready_o         (ready_60_to_50_v0),
    .vert0_data_o          (data_60_to_70_v0),
    .vert0_valid_o         (valid_60_to_70_v0),
    .vert0_ready_i         (ready_70_to_60_v0),
    .vert1_data_i          (data_50_to_60_v1),
    .vert1_valid_i         (valid_50_to_60_v1),
    .vert1_ready_o         (ready_60_to_50_v1),
    .vert1_data_o          (data_60_to_70_v1),
    .vert1_valid_o         (valid_60_to_70_v1),
    .vert1_ready_i         (ready_70_to_60_v1),
    .local_data_i          (data_i[0][6]),
    .local_valid_i         (valid_i[0][6]),
    .local_ready_o         (ready_o[0][6]),
    .local_data_o          (data_o[0][6]),
    .local_valid_o         (valid_o[0][6]),
    .local_ready_i         (ready_i[0][6]),
    .credit_upd            (credit_upd)
);

/*Router 0,7*/    
cast_router #(
    .isUBM_list            (isUBM_list_0_7),
    .isFC_list             (isFC_list_0_7),
    .FCdn_list             (FCdn_list_0_7),
    .FCpl_list             (FCpl_list_0_7),
    .rt_file_list          (cast_rt_file_list_0_7)
)router_0_7(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (34'b0),
    .west_valid_i          (1'b0),
    .west_ready_o          (),
    .west_data_o           (),
    .west_valid_o          (),
    .west_ready_i          (1'b0),
    .east_data_i           (data_71_to_70),
    .east_valid_i          (valid_71_to_70),
    .east_ready_o          (ready_70_to_71),
    .east_data_o           (data_70_to_71),
    .east_valid_o          (valid_70_to_71),
    .east_ready_i          (ready_71_to_70),
    .vert0_data_i          (data_60_to_70_v0),
    .vert0_valid_i         (valid_60_to_70_v0),
    .vert0_ready_o         (ready_70_to_60_v0),
    .vert0_data_o          (data_70_to_80_v0),
    .vert0_valid_o         (valid_70_to_80_v0),
    .vert0_ready_i         (ready_80_to_70_v0),
    .vert1_data_i          (data_60_to_70_v1),
    .vert1_valid_i         (valid_60_to_70_v1),
    .vert1_ready_o         (ready_70_to_60_v1),
    .vert1_data_o          (data_70_to_80_v1),
    .vert1_valid_o         (valid_70_to_80_v1),
    .vert1_ready_i         (ready_80_to_70_v1),
    .local_data_i          (data_i[0][7]),
    .local_valid_i         (valid_i[0][7]),
    .local_ready_o         (ready_o[0][7]),
    .local_data_o          (data_o[0][7]),
    .local_valid_o         (valid_o[0][7]),
    .local_ready_i         (ready_i[0][7]),
    .credit_upd            (credit_upd)
);

/*Router 0,8*/    
cast_router #(
    .isUBM_list            (isUBM_list_0_8),
    .isFC_list             (isFC_list_0_8),
    .FCdn_list             (FCdn_list_0_8),
    .FCpl_list             (FCpl_list_0_8),
    .rt_file_list          (cast_rt_file_list_0_8)
)router_0_8(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (34'b0),
    .west_valid_i          (1'b0),
    .west_ready_o          (),
    .west_data_o           (),
    .west_valid_o          (),
    .west_ready_i          (1'b0),
    .east_data_i           (data_81_to_80),
    .east_valid_i          (valid_81_to_80),
    .east_ready_o          (ready_80_to_81),
    .east_data_o           (data_80_to_81),
    .east_valid_o          (valid_80_to_81),
    .east_ready_i          (ready_81_to_80),
    .vert0_data_i          (data_70_to_80_v0),
    .vert0_valid_i         (valid_70_to_80_v0),
    .vert0_ready_o         (ready_80_to_70_v0),
    .vert0_data_o          (data_80_to_90_v0),
    .vert0_valid_o         (valid_80_to_90_v0),
    .vert0_ready_i         (ready_90_to_80_v0),
    .vert1_data_i          (data_70_to_80_v1),
    .vert1_valid_i         (valid_70_to_80_v1),
    .vert1_ready_o         (ready_80_to_70_v1),
    .vert1_data_o          (data_80_to_90_v1),
    .vert1_valid_o         (valid_80_to_90_v1),
    .vert1_ready_i         (ready_90_to_80_v1),
    .local_data_i          (data_i[0][8]),
    .local_valid_i         (valid_i[0][8]),
    .local_ready_o         (ready_o[0][8]),
    .local_data_o          (data_o[0][8]),
    .local_valid_o         (valid_o[0][8]),
    .local_ready_i         (ready_i[0][8]),
    .credit_upd            (credit_upd)
);

/*Router 0,9*/    
cast_router #(
    .isUBM_list            (isUBM_list_0_9),
    .isFC_list             (isFC_list_0_9),
    .FCdn_list             (FCdn_list_0_9),
    .FCpl_list             (FCpl_list_0_9),
    .rt_file_list          (cast_rt_file_list_0_9)
)router_0_9(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (34'b0),
    .west_valid_i          (1'b0),
    .west_ready_o          (),
    .west_data_o           (),
    .west_valid_o          (),
    .west_ready_i          (1'b0),
    .east_data_i           (data_91_to_90),
    .east_valid_i          (valid_91_to_90),
    .east_ready_o          (ready_90_to_91),
    .east_data_o           (data_90_to_91),
    .east_valid_o          (valid_90_to_91),
    .east_ready_i          (ready_91_to_90),
    .vert0_data_i          (data_80_to_90_v0),
    .vert0_valid_i         (valid_80_to_90_v0),
    .vert0_ready_o         (ready_90_to_80_v0),
    .vert0_data_o          (data_90_to_100_v0),
    .vert0_valid_o         (valid_90_to_100_v0),
    .vert0_ready_i         (ready_100_to_90_v0),
    .vert1_data_i          (data_80_to_90_v1),
    .vert1_valid_i         (valid_80_to_90_v1),
    .vert1_ready_o         (ready_90_to_80_v1),
    .vert1_data_o          (data_90_to_100_v1),
    .vert1_valid_o         (valid_90_to_100_v1),
    .vert1_ready_i         (ready_100_to_90_v1),
    .local_data_i          (data_i[0][9]),
    .local_valid_i         (valid_i[0][9]),
    .local_ready_o         (ready_o[0][9]),
    .local_data_o          (data_o[0][9]),
    .local_valid_o         (valid_o[0][9]),
    .local_ready_i         (ready_i[0][9]),
    .credit_upd            (credit_upd)
);

/*Router 0,10*/    
cast_router #(
    .isUBM_list            (isUBM_list_0_10),
    .isFC_list             (isFC_list_0_10),
    .FCdn_list             (FCdn_list_0_10),
    .FCpl_list             (FCpl_list_0_10),
    .rt_file_list          (cast_rt_file_list_0_10)
)router_0_10(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (34'b0),
    .west_valid_i          (1'b0),
    .west_ready_o          (),
    .west_data_o           (),
    .west_valid_o          (),
    .west_ready_i          (1'b0),
    .east_data_i           (data_101_to_100),
    .east_valid_i          (valid_101_to_100),
    .east_ready_o          (ready_100_to_101),
    .east_data_o           (data_100_to_101),
    .east_valid_o          (valid_100_to_101),
    .east_ready_i          (ready_101_to_100),
    .vert0_data_i          (data_90_to_100_v0),
    .vert0_valid_i         (valid_90_to_100_v0),
    .vert0_ready_o         (ready_100_to_90_v0),
    .vert0_data_o          (data_100_to_110_v0),
    .vert0_valid_o         (valid_100_to_110_v0),
    .vert0_ready_i         (ready_110_to_100_v0),
    .vert1_data_i          (data_90_to_100_v1),
    .vert1_valid_i         (valid_90_to_100_v1),
    .vert1_ready_o         (ready_100_to_90_v1),
    .vert1_data_o          (data_100_to_110_v1),
    .vert1_valid_o         (valid_100_to_110_v1),
    .vert1_ready_i         (ready_110_to_100_v1),
    .local_data_i          (data_i[0][10]),
    .local_valid_i         (valid_i[0][10]),
    .local_ready_o         (ready_o[0][10]),
    .local_data_o          (data_o[0][10]),
    .local_valid_o         (valid_o[0][10]),
    .local_ready_i         (ready_i[0][10]),
    .credit_upd            (credit_upd)
);

/*Router 0,11*/    
cast_router #(
    .isUBM_list            (isUBM_list_0_11),
    .isFC_list             (isFC_list_0_11),
    .FCdn_list             (FCdn_list_0_11),
    .FCpl_list             (FCpl_list_0_11),
    .rt_file_list          (cast_rt_file_list_0_11)
)router_0_11(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (34'b0),
    .west_valid_i          (1'b0),
    .west_ready_o          (),
    .west_data_o           (),
    .west_valid_o          (),
    .west_ready_i          (1'b0),
    .east_data_i           (data_111_to_110),
    .east_valid_i          (valid_111_to_110),
    .east_ready_o          (ready_110_to_111),
    .east_data_o           (data_110_to_111),
    .east_valid_o          (valid_110_to_111),
    .east_ready_i          (ready_111_to_110),
    .vert0_data_i          (data_100_to_110_v0),
    .vert0_valid_i         (valid_100_to_110_v0),
    .vert0_ready_o         (ready_110_to_100_v0),
    .vert0_data_o          (data_110_to_120_v0),
    .vert0_valid_o         (valid_110_to_120_v0),
    .vert0_ready_i         (ready_120_to_110_v0),
    .vert1_data_i          (data_100_to_110_v1),
    .vert1_valid_i         (valid_100_to_110_v1),
    .vert1_ready_o         (ready_110_to_100_v1),
    .vert1_data_o          (data_110_to_120_v1),
    .vert1_valid_o         (valid_110_to_120_v1),
    .vert1_ready_i         (ready_120_to_110_v1),
    .local_data_i          (data_i[0][11]),
    .local_valid_i         (valid_i[0][11]),
    .local_ready_o         (ready_o[0][11]),
    .local_data_o          (data_o[0][11]),
    .local_valid_o         (valid_o[0][11]),
    .local_ready_i         (ready_i[0][11]),
    .credit_upd            (credit_upd)
);

/*Router 0,12*/    
cast_router #(
    .isUBM_list            (isUBM_list_0_12),
    .isFC_list             (isFC_list_0_12),
    .FCdn_list             (FCdn_list_0_12),
    .FCpl_list             (FCpl_list_0_12),
    .rt_file_list          (cast_rt_file_list_0_12)
)router_0_12(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (34'b0),
    .west_valid_i          (1'b0),
    .west_ready_o          (),
    .west_data_o           (),
    .west_valid_o          (),
    .west_ready_i          (1'b0),
    .east_data_i           (data_121_to_120),
    .east_valid_i          (valid_121_to_120),
    .east_ready_o          (ready_120_to_121),
    .east_data_o           (data_120_to_121),
    .east_valid_o          (valid_120_to_121),
    .east_ready_i          (ready_121_to_120),
    .vert0_data_i          (data_110_to_120_v0),
    .vert0_valid_i         (valid_110_to_120_v0),
    .vert0_ready_o         (ready_120_to_110_v0),
    .vert0_data_o          (data_120_to_130_v0),
    .vert0_valid_o         (valid_120_to_130_v0),
    .vert0_ready_i         (ready_130_to_120_v0),
    .vert1_data_i          (data_110_to_120_v1),
    .vert1_valid_i         (valid_110_to_120_v1),
    .vert1_ready_o         (ready_120_to_110_v1),
    .vert1_data_o          (data_120_to_130_v1),
    .vert1_valid_o         (valid_120_to_130_v1),
    .vert1_ready_i         (ready_130_to_120_v1),
    .local_data_i          (data_i[0][12]),
    .local_valid_i         (valid_i[0][12]),
    .local_ready_o         (ready_o[0][12]),
    .local_data_o          (data_o[0][12]),
    .local_valid_o         (valid_o[0][12]),
    .local_ready_i         (ready_i[0][12]),
    .credit_upd            (credit_upd)
);

/*Router 0,13*/    
cast_router #(
    .isUBM_list            (isUBM_list_0_13),
    .isFC_list             (isFC_list_0_13),
    .FCdn_list             (FCdn_list_0_13),
    .FCpl_list             (FCpl_list_0_13),
    .rt_file_list          (cast_rt_file_list_0_13)
)router_0_13(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (34'b0),
    .west_valid_i          (1'b0),
    .west_ready_o          (),
    .west_data_o           (),
    .west_valid_o          (),
    .west_ready_i          (1'b0),
    .east_data_i           (data_131_to_130),
    .east_valid_i          (valid_131_to_130),
    .east_ready_o          (ready_130_to_131),
    .east_data_o           (data_130_to_131),
    .east_valid_o          (valid_130_to_131),
    .east_ready_i          (ready_131_to_130),
    .vert0_data_i          (data_120_to_130_v0),
    .vert0_valid_i         (valid_120_to_130_v0),
    .vert0_ready_o         (ready_130_to_120_v0),
    .vert0_data_o          (data_130_to_140_v0),
    .vert0_valid_o         (valid_130_to_140_v0),
    .vert0_ready_i         (ready_140_to_130_v0),
    .vert1_data_i          (data_120_to_130_v1),
    .vert1_valid_i         (valid_120_to_130_v1),
    .vert1_ready_o         (ready_130_to_120_v1),
    .vert1_data_o          (data_130_to_140_v1),
    .vert1_valid_o         (valid_130_to_140_v1),
    .vert1_ready_i         (ready_140_to_130_v1),
    .local_data_i          (data_i[0][13]),
    .local_valid_i         (valid_i[0][13]),
    .local_ready_o         (ready_o[0][13]),
    .local_data_o          (data_o[0][13]),
    .local_valid_o         (valid_o[0][13]),
    .local_ready_i         (ready_i[0][13]),
    .credit_upd            (credit_upd)
);

/*Router 0,14*/    
cast_router #(
    .isUBM_list            (isUBM_list_0_14),
    .isFC_list             (isFC_list_0_14),
    .FCdn_list             (FCdn_list_0_14),
    .FCpl_list             (FCpl_list_0_14),
    .rt_file_list          (cast_rt_file_list_0_14)
)router_0_14(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (34'b0),
    .west_valid_i          (1'b0),
    .west_ready_o          (),
    .west_data_o           (),
    .west_valid_o          (),
    .west_ready_i          (1'b0),
    .east_data_i           (data_141_to_140),
    .east_valid_i          (valid_141_to_140),
    .east_ready_o          (ready_140_to_141),
    .east_data_o           (data_140_to_141),
    .east_valid_o          (valid_140_to_141),
    .east_ready_i          (ready_141_to_140),
    .vert0_data_i          (data_130_to_140_v0),
    .vert0_valid_i         (valid_130_to_140_v0),
    .vert0_ready_o         (ready_140_to_130_v0),
    .vert0_data_o          (data_140_to_150_v0),
    .vert0_valid_o         (valid_140_to_150_v0),
    .vert0_ready_i         (ready_150_to_140_v0),
    .vert1_data_i          (data_130_to_140_v1),
    .vert1_valid_i         (valid_130_to_140_v1),
    .vert1_ready_o         (ready_140_to_130_v1),
    .vert1_data_o          (data_140_to_150_v1),
    .vert1_valid_o         (valid_140_to_150_v1),
    .vert1_ready_i         (ready_150_to_140_v1),
    .local_data_i          (data_i[0][14]),
    .local_valid_i         (valid_i[0][14]),
    .local_ready_o         (ready_o[0][14]),
    .local_data_o          (data_o[0][14]),
    .local_valid_o         (valid_o[0][14]),
    .local_ready_i         (ready_i[0][14]),
    .credit_upd            (credit_upd)
);

/*Router 0,15*/    
cast_router #(
    .isUBM_list            (isUBM_list_0_15),
    .isFC_list             (isFC_list_0_15),
    .FCdn_list             (FCdn_list_0_15),
    .FCpl_list             (FCpl_list_0_15),
    .rt_file_list          (cast_rt_file_list_0_15)
)router_0_15(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (34'b0),
    .west_valid_i          (1'b0),
    .west_ready_o          (),
    .west_data_o           (),
    .west_valid_o          (),
    .west_ready_i          (1'b0),
    .east_data_i           (data_151_to_150),
    .east_valid_i          (valid_151_to_150),
    .east_ready_o          (ready_150_to_151),
    .east_data_o           (data_150_to_151),
    .east_valid_o          (valid_150_to_151),
    .east_ready_i          (ready_151_to_150),
    .vert0_data_i          (data_140_to_150_v0),
    .vert0_valid_i         (valid_140_to_150_v0),
    .vert0_ready_o         (ready_150_to_140_v0),
    .vert0_data_o          (data_150_to_160_v0),
    .vert0_valid_o         (valid_150_to_160_v0),
    .vert0_ready_i         (ready_160_to_150_v0),
    .vert1_data_i          (data_140_to_150_v1),
    .vert1_valid_i         (valid_140_to_150_v1),
    .vert1_ready_o         (ready_150_to_140_v1),
    .vert1_data_o          (data_150_to_160_v1),
    .vert1_valid_o         (valid_150_to_160_v1),
    .vert1_ready_i         (ready_160_to_150_v1),
    .local_data_i          (data_i[0][15]),
    .local_valid_i         (valid_i[0][15]),
    .local_ready_o         (ready_o[0][15]),
    .local_data_o          (data_o[0][15]),
    .local_valid_o         (valid_o[0][15]),
    .local_ready_i         (ready_i[0][15]),
    .credit_upd            (credit_upd)
);

/*Router 0,16*/    
cast_router #(
    .isUBM_list            (isUBM_list_0_16),
    .isFC_list             (isFC_list_0_16),
    .FCdn_list             (FCdn_list_0_16),
    .FCpl_list             (FCpl_list_0_16),
    .rt_file_list          (cast_rt_file_list_0_16)
)router_0_16(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (34'b0),
    .west_valid_i          (1'b0),
    .west_ready_o          (),
    .west_data_o           (),
    .west_valid_o          (),
    .west_ready_i          (1'b0),
    .east_data_i           (data_161_to_160),
    .east_valid_i          (valid_161_to_160),
    .east_ready_o          (ready_160_to_161),
    .east_data_o           (data_160_to_161),
    .east_valid_o          (valid_160_to_161),
    .east_ready_i          (ready_161_to_160),
    .vert0_data_i          (data_150_to_160_v0),
    .vert0_valid_i         (valid_150_to_160_v0),
    .vert0_ready_o         (ready_160_to_150_v0),
    .vert0_data_o          (data_160_to_170_v0),
    .vert0_valid_o         (valid_160_to_170_v0),
    .vert0_ready_i         (ready_170_to_160_v0),
    .vert1_data_i          (data_150_to_160_v1),
    .vert1_valid_i         (valid_150_to_160_v1),
    .vert1_ready_o         (ready_160_to_150_v1),
    .vert1_data_o          (data_160_to_170_v1),
    .vert1_valid_o         (valid_160_to_170_v1),
    .vert1_ready_i         (ready_170_to_160_v1),
    .local_data_i          (data_i[0][16]),
    .local_valid_i         (valid_i[0][16]),
    .local_ready_o         (ready_o[0][16]),
    .local_data_o          (data_o[0][16]),
    .local_valid_o         (valid_o[0][16]),
    .local_ready_i         (ready_i[0][16]),
    .credit_upd            (credit_upd)
);

/*Router 0,17*/    
cast_router #(
    .isUBM_list            (isUBM_list_0_17),
    .isFC_list             (isFC_list_0_17),
    .FCdn_list             (FCdn_list_0_17),
    .FCpl_list             (FCpl_list_0_17),
    .rt_file_list          (cast_rt_file_list_0_17)
)router_0_17(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (34'b0),
    .west_valid_i          (1'b0),
    .west_ready_o          (),
    .west_data_o           (),
    .west_valid_o          (),
    .west_ready_i          (1'b0),
    .east_data_i           (data_171_to_170),
    .east_valid_i          (valid_171_to_170),
    .east_ready_o          (ready_170_to_171),
    .east_data_o           (data_170_to_171),
    .east_valid_o          (valid_170_to_171),
    .east_ready_i          (ready_171_to_170),
    .vert0_data_i          (data_160_to_170_v0),
    .vert0_valid_i         (valid_160_to_170_v0),
    .vert0_ready_o         (ready_170_to_160_v0),
    .vert0_data_o          (data_170_to_180_v0),
    .vert0_valid_o         (valid_170_to_180_v0),
    .vert0_ready_i         (ready_180_to_170_v0),
    .vert1_data_i          (data_160_to_170_v1),
    .vert1_valid_i         (valid_160_to_170_v1),
    .vert1_ready_o         (ready_170_to_160_v1),
    .vert1_data_o          (data_170_to_180_v1),
    .vert1_valid_o         (valid_170_to_180_v1),
    .vert1_ready_i         (ready_180_to_170_v1),
    .local_data_i          (data_i[0][17]),
    .local_valid_i         (valid_i[0][17]),
    .local_ready_o         (ready_o[0][17]),
    .local_data_o          (data_o[0][17]),
    .local_valid_o         (valid_o[0][17]),
    .local_ready_i         (ready_i[0][17]),
    .credit_upd            (credit_upd)
);

/*Router 0,18*/    
cast_router #(
    .isUBM_list            (isUBM_list_0_18),
    .isFC_list             (isFC_list_0_18),
    .FCdn_list             (FCdn_list_0_18),
    .FCpl_list             (FCpl_list_0_18),
    .rt_file_list          (cast_rt_file_list_0_18)
)router_0_18(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (34'b0),
    .west_valid_i          (1'b0),
    .west_ready_o          (),
    .west_data_o           (),
    .west_valid_o          (),
    .west_ready_i          (1'b0),
    .east_data_i           (data_181_to_180),
    .east_valid_i          (valid_181_to_180),
    .east_ready_o          (ready_180_to_181),
    .east_data_o           (data_180_to_181),
    .east_valid_o          (valid_180_to_181),
    .east_ready_i          (ready_181_to_180),
    .vert0_data_i          (data_170_to_180_v0),
    .vert0_valid_i         (valid_170_to_180_v0),
    .vert0_ready_o         (ready_180_to_170_v0),
    .vert0_data_o          (data_180_to_190_v0),
    .vert0_valid_o         (valid_180_to_190_v0),
    .vert0_ready_i         (ready_190_to_180_v0),
    .vert1_data_i          (data_170_to_180_v1),
    .vert1_valid_i         (valid_170_to_180_v1),
    .vert1_ready_o         (ready_180_to_170_v1),
    .vert1_data_o          (data_180_to_190_v1),
    .vert1_valid_o         (valid_180_to_190_v1),
    .vert1_ready_i         (ready_190_to_180_v1),
    .local_data_i          (data_i[0][18]),
    .local_valid_i         (valid_i[0][18]),
    .local_ready_o         (ready_o[0][18]),
    .local_data_o          (data_o[0][18]),
    .local_valid_o         (valid_o[0][18]),
    .local_ready_i         (ready_i[0][18]),
    .credit_upd            (credit_upd)
);

/*Router 0,19*/    
cast_router #(
    .isUBM_list            (isUBM_list_0_19),
    .isFC_list             (isFC_list_0_19),
    .FCdn_list             (FCdn_list_0_19),
    .FCpl_list             (FCpl_list_0_19),
    .rt_file_list          (cast_rt_file_list_0_19)
)router_0_19(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (34'b0),
    .west_valid_i          (1'b0),
    .west_ready_o          (),
    .west_data_o           (),
    .west_valid_o          (),
    .west_ready_i          (1'b0),
    .east_data_i           (data_191_to_190),
    .east_valid_i          (valid_191_to_190),
    .east_ready_o          (ready_190_to_191),
    .east_data_o           (data_190_to_191),
    .east_valid_o          (valid_190_to_191),
    .east_ready_i          (ready_191_to_190),
    .vert0_data_i          (data_180_to_190_v0),
    .vert0_valid_i         (valid_180_to_190_v0),
    .vert0_ready_o         (ready_190_to_180_v0),
    .vert0_data_o          (data_190_to_200_v0),
    .vert0_valid_o         (valid_190_to_200_v0),
    .vert0_ready_i         (ready_200_to_190_v0),
    .vert1_data_i          (data_180_to_190_v1),
    .vert1_valid_i         (valid_180_to_190_v1),
    .vert1_ready_o         (ready_190_to_180_v1),
    .vert1_data_o          (data_190_to_200_v1),
    .vert1_valid_o         (valid_190_to_200_v1),
    .vert1_ready_i         (ready_200_to_190_v1),
    .local_data_i          (data_i[0][19]),
    .local_valid_i         (valid_i[0][19]),
    .local_ready_o         (ready_o[0][19]),
    .local_data_o          (data_o[0][19]),
    .local_valid_o         (valid_o[0][19]),
    .local_ready_i         (ready_i[0][19]),
    .credit_upd            (credit_upd)
);

/*Router 0,20*/    
cast_router #(
    .isUBM_list            (isUBM_list_0_20),
    .isFC_list             (isFC_list_0_20),
    .FCdn_list             (FCdn_list_0_20),
    .FCpl_list             (FCpl_list_0_20),
    .rt_file_list          (cast_rt_file_list_0_20)
)router_0_20(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (34'b0),
    .west_valid_i          (1'b0),
    .west_ready_o          (),
    .west_data_o           (),
    .west_valid_o          (),
    .west_ready_i          (1'b0),
    .east_data_i           (data_201_to_200),
    .east_valid_i          (valid_201_to_200),
    .east_ready_o          (ready_200_to_201),
    .east_data_o           (data_200_to_201),
    .east_valid_o          (valid_200_to_201),
    .east_ready_i          (ready_201_to_200),
    .vert0_data_i          (data_190_to_200_v0),
    .vert0_valid_i         (valid_190_to_200_v0),
    .vert0_ready_o         (ready_200_to_190_v0),
    .vert0_data_o          (data_200_to_210_v0),
    .vert0_valid_o         (valid_200_to_210_v0),
    .vert0_ready_i         (ready_210_to_200_v0),
    .vert1_data_i          (data_190_to_200_v1),
    .vert1_valid_i         (valid_190_to_200_v1),
    .vert1_ready_o         (ready_200_to_190_v1),
    .vert1_data_o          (data_200_to_210_v1),
    .vert1_valid_o         (valid_200_to_210_v1),
    .vert1_ready_i         (ready_210_to_200_v1),
    .local_data_i          (data_i[0][20]),
    .local_valid_i         (valid_i[0][20]),
    .local_ready_o         (ready_o[0][20]),
    .local_data_o          (data_o[0][20]),
    .local_valid_o         (valid_o[0][20]),
    .local_ready_i         (ready_i[0][20]),
    .credit_upd            (credit_upd)
);

/*Router 0,21*/    
cast_router #(
    .isUBM_list            (isUBM_list_0_21),
    .isFC_list             (isFC_list_0_21),
    .FCdn_list             (FCdn_list_0_21),
    .FCpl_list             (FCpl_list_0_21),
    .rt_file_list          (cast_rt_file_list_0_21)
)router_0_21(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (34'b0),
    .west_valid_i          (1'b0),
    .west_ready_o          (),
    .west_data_o           (),
    .west_valid_o          (),
    .west_ready_i          (1'b0),
    .east_data_i           (data_211_to_210),
    .east_valid_i          (valid_211_to_210),
    .east_ready_o          (ready_210_to_211),
    .east_data_o           (data_210_to_211),
    .east_valid_o          (valid_210_to_211),
    .east_ready_i          (ready_211_to_210),
    .vert0_data_i          (data_200_to_210_v0),
    .vert0_valid_i         (valid_200_to_210_v0),
    .vert0_ready_o         (ready_210_to_200_v0),
    .vert0_data_o          (data_210_to_220_v0),
    .vert0_valid_o         (valid_210_to_220_v0),
    .vert0_ready_i         (ready_220_to_210_v0),
    .vert1_data_i          (data_200_to_210_v1),
    .vert1_valid_i         (valid_200_to_210_v1),
    .vert1_ready_o         (ready_210_to_200_v1),
    .vert1_data_o          (data_210_to_220_v1),
    .vert1_valid_o         (valid_210_to_220_v1),
    .vert1_ready_i         (ready_220_to_210_v1),
    .local_data_i          (data_i[0][21]),
    .local_valid_i         (valid_i[0][21]),
    .local_ready_o         (ready_o[0][21]),
    .local_data_o          (data_o[0][21]),
    .local_valid_o         (valid_o[0][21]),
    .local_ready_i         (ready_i[0][21]),
    .credit_upd            (credit_upd)
);

/*Router 0,22*/    
cast_router #(
    .isUBM_list            (isUBM_list_0_22),
    .isFC_list             (isFC_list_0_22),
    .FCdn_list             (FCdn_list_0_22),
    .FCpl_list             (FCpl_list_0_22),
    .rt_file_list          (cast_rt_file_list_0_22)
)router_0_22(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (34'b0),
    .west_valid_i          (1'b0),
    .west_ready_o          (),
    .west_data_o           (),
    .west_valid_o          (),
    .west_ready_i          (1'b0),
    .east_data_i           (data_221_to_220),
    .east_valid_i          (valid_221_to_220),
    .east_ready_o          (ready_220_to_221),
    .east_data_o           (data_220_to_221),
    .east_valid_o          (valid_220_to_221),
    .east_ready_i          (ready_221_to_220),
    .vert0_data_i          (data_210_to_220_v0),
    .vert0_valid_i         (valid_210_to_220_v0),
    .vert0_ready_o         (ready_220_to_210_v0),
    .vert0_data_o          (data_220_to_230_v0),
    .vert0_valid_o         (valid_220_to_230_v0),
    .vert0_ready_i         (ready_230_to_220_v0),
    .vert1_data_i          (data_210_to_220_v1),
    .vert1_valid_i         (valid_210_to_220_v1),
    .vert1_ready_o         (ready_220_to_210_v1),
    .vert1_data_o          (data_220_to_230_v1),
    .vert1_valid_o         (valid_220_to_230_v1),
    .vert1_ready_i         (ready_230_to_220_v1),
    .local_data_i          (data_i[0][22]),
    .local_valid_i         (valid_i[0][22]),
    .local_ready_o         (ready_o[0][22]),
    .local_data_o          (data_o[0][22]),
    .local_valid_o         (valid_o[0][22]),
    .local_ready_i         (ready_i[0][22]),
    .credit_upd            (credit_upd)
);

/*Router 0,23*/    
cast_router #(
    .isUBM_list            (isUBM_list_0_23),
    .isFC_list             (isFC_list_0_23),
    .FCdn_list             (FCdn_list_0_23),
    .FCpl_list             (FCpl_list_0_23),
    .rt_file_list          (cast_rt_file_list_0_23)
)router_0_23(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (34'b0),
    .west_valid_i          (1'b0),
    .west_ready_o          (),
    .west_data_o           (data_o_flee6),
    .west_valid_o          (valid_o_flee6),
    .west_ready_i          (ready_i_flee6),
    .east_data_i           (data_231_to_230),
    .east_valid_i          (valid_231_to_230),
    .east_ready_o          (ready_230_to_231),
    .east_data_o           (data_230_to_231),
    .east_valid_o          (valid_230_to_231),
    .east_ready_i          (ready_231_to_230),
    .vert0_data_i          (data_220_to_230_v0),
    .vert0_valid_i         (valid_220_to_230_v0),
    .vert0_ready_o         (ready_230_to_220_v0),
    .vert0_data_o          (data_230_to_240_v0),
    .vert0_valid_o         (valid_230_to_240_v0),
    .vert0_ready_i         (ready_240_to_230_v0),
    .vert1_data_i          (data_220_to_230_v1),
    .vert1_valid_i         (valid_220_to_230_v1),
    .vert1_ready_o         (ready_230_to_220_v1),
    .vert1_data_o          (data_230_to_240_v1),
    .vert1_valid_o         (valid_230_to_240_v1),
    .vert1_ready_i         (ready_240_to_230_v1),
    .local_data_i          (data_i[0][23]),
    .local_valid_i         (valid_i[0][23]),
    .local_ready_o         (ready_o[0][23]),
    .local_data_o          (data_o[0][23]),
    .local_valid_o         (valid_o[0][23]),
    .local_ready_i         (ready_i[0][23]),
    .credit_upd            (credit_upd)
);

/*Router 0,24*/    
cast_router #(
    .isUBM_list            (isUBM_list_0_24),
    .isFC_list             (isFC_list_0_24),
    .FCdn_list             (FCdn_list_0_24),
    .FCpl_list             (FCpl_list_0_24),
    .rt_file_list          (cast_rt_file_list_0_24)
)router_0_24(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (34'b0),
    .west_valid_i          (1'b0),
    .west_ready_o          (),
    .west_data_o           (),
    .west_valid_o          (),
    .west_ready_i          (1'b0),
    .east_data_i           (data_241_to_240),
    .east_valid_i          (valid_241_to_240),
    .east_ready_o          (ready_240_to_241),
    .east_data_o           (data_240_to_241),
    .east_valid_o          (valid_240_to_241),
    .east_ready_i          (ready_241_to_240),
    .vert0_data_i          (data_230_to_240_v0),
    .vert0_valid_i         (valid_230_to_240_v0),
    .vert0_ready_o         (ready_240_to_230_v0),
    .vert0_data_o          (),
    .vert0_valid_o         (),
    .vert0_ready_i         (1'b0),
    .vert1_data_i          (data_230_to_240_v1),
    .vert1_valid_i         (valid_230_to_240_v1),
    .vert1_ready_o         (ready_240_to_230_v1),
    .vert1_data_o          (),
    .vert1_valid_o         (),
    .vert1_ready_i         (1'b0),
    .local_data_i          (data_i[0][24]),
    .local_valid_i         (valid_i[0][24]),
    .local_ready_o         (ready_o[0][24]),
    .local_data_o          (data_o[0][24]),
    .local_valid_o         (valid_o[0][24]),
    .local_ready_i         (ready_i[0][24]),
    .credit_upd            (credit_upd)
);

/*Router 1,0*/    
cast_router #(
    .isUBM_list            (isUBM_list_1_0),
    .isFC_list             (isFC_list_1_0),
    .FCdn_list             (FCdn_list_1_0),
    .FCpl_list             (FCpl_list_1_0),
    .rt_file_list          (cast_rt_file_list_1_0)
)router_1_0(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_0_to_1),
    .west_valid_i          (valid_0_to_1),
    .west_ready_o          (ready_1_to_0),
    .west_data_o           (data_1_to_0),
    .west_valid_o          (valid_1_to_0),
    .west_ready_i          (ready_0_to_1),
    .east_data_i           (data_2_to_1),
    .east_valid_i          (valid_2_to_1),
    .east_ready_o          (ready_1_to_2),
    .east_data_o           (data_1_to_2),
    .east_valid_o          (valid_1_to_2),
    .east_ready_i          (ready_2_to_1),
    .vert0_data_i          (34'b0),
    .vert0_valid_i         (1'b0),
    .vert0_ready_o         (),
    .vert0_data_o          (data_1_to_11_v0),
    .vert0_valid_o         (valid_1_to_11_v0),
    .vert0_ready_i         (ready_11_to_1_v0),
    .vert1_data_i          (34'b0),
    .vert1_valid_i         (1'b0),
    .vert1_ready_o         (),
    .vert1_data_o          (data_1_to_11_v1),
    .vert1_valid_o         (valid_1_to_11_v1),
    .vert1_ready_i         (ready_11_to_1_v1),
    .local_data_i          (data_i[1][0]),
    .local_valid_i         (valid_i[1][0]),
    .local_ready_o         (ready_o[1][0]),
    .local_data_o          (data_o[1][0]),
    .local_valid_o         (valid_o[1][0]),
    .local_ready_i         (ready_i[1][0]),
    .credit_upd            (credit_upd)
);

/*Router 1,1*/    
cast_router #(
    .isUBM_list            (isUBM_list_1_1),
    .isFC_list             (isFC_list_1_1),
    .FCdn_list             (FCdn_list_1_1),
    .FCpl_list             (FCpl_list_1_1),
    .rt_file_list          (cast_rt_file_list_1_1)
)router_1_1(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_10_to_11),
    .west_valid_i          (valid_10_to_11),
    .west_ready_o          (ready_11_to_10),
    .west_data_o           (data_11_to_10),
    .west_valid_o          (valid_11_to_10),
    .west_ready_i          (ready_10_to_11),
    .east_data_i           (data_12_to_11),
    .east_valid_i          (valid_12_to_11),
    .east_ready_o          (ready_11_to_12),
    .east_data_o           (data_11_to_12),
    .east_valid_o          (valid_11_to_12),
    .east_ready_i          (ready_12_to_11),
    .vert0_data_i          (data_1_to_11_v0),
    .vert0_valid_i         (valid_1_to_11_v0),
    .vert0_ready_o         (ready_11_to_1_v0),
    .vert0_data_o          (data_11_to_21_v0),
    .vert0_valid_o         (valid_11_to_21_v0),
    .vert0_ready_i         (ready_21_to_11_v0),
    .vert1_data_i          (data_1_to_11_v1),
    .vert1_valid_i         (valid_1_to_11_v1),
    .vert1_ready_o         (ready_11_to_1_v1),
    .vert1_data_o          (data_11_to_21_v1),
    .vert1_valid_o         (valid_11_to_21_v1),
    .vert1_ready_i         (ready_21_to_11_v1),
    .local_data_i          (data_i[1][1]),
    .local_valid_i         (valid_i[1][1]),
    .local_ready_o         (ready_o[1][1]),
    .local_data_o          (data_o[1][1]),
    .local_valid_o         (valid_o[1][1]),
    .local_ready_i         (ready_i[1][1]),
    .credit_upd            (credit_upd)
);

/*Router 1,2*/    
cast_router #(
    .isUBM_list            (isUBM_list_1_2),
    .isFC_list             (isFC_list_1_2),
    .FCdn_list             (FCdn_list_1_2),
    .FCpl_list             (FCpl_list_1_2),
    .rt_file_list          (cast_rt_file_list_1_2)
)router_1_2(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_20_to_21),
    .west_valid_i          (valid_20_to_21),
    .west_ready_o          (ready_21_to_20),
    .west_data_o           (data_21_to_20),
    .west_valid_o          (valid_21_to_20),
    .west_ready_i          (ready_20_to_21),
    .east_data_i           (data_22_to_21),
    .east_valid_i          (valid_22_to_21),
    .east_ready_o          (ready_21_to_22),
    .east_data_o           (data_21_to_22),
    .east_valid_o          (valid_21_to_22),
    .east_ready_i          (ready_22_to_21),
    .vert0_data_i          (data_11_to_21_v0),
    .vert0_valid_i         (valid_11_to_21_v0),
    .vert0_ready_o         (ready_21_to_11_v0),
    .vert0_data_o          (data_21_to_31_v0),
    .vert0_valid_o         (valid_21_to_31_v0),
    .vert0_ready_i         (ready_31_to_21_v0),
    .vert1_data_i          (data_11_to_21_v1),
    .vert1_valid_i         (valid_11_to_21_v1),
    .vert1_ready_o         (ready_21_to_11_v1),
    .vert1_data_o          (data_21_to_31_v1),
    .vert1_valid_o         (valid_21_to_31_v1),
    .vert1_ready_i         (ready_31_to_21_v1),
    .local_data_i          (data_i[1][2]),
    .local_valid_i         (valid_i[1][2]),
    .local_ready_o         (ready_o[1][2]),
    .local_data_o          (data_o[1][2]),
    .local_valid_o         (valid_o[1][2]),
    .local_ready_i         (ready_i[1][2]),
    .credit_upd            (credit_upd)
);

/*Router 1,3*/    
cast_router #(
    .isUBM_list            (isUBM_list_1_3),
    .isFC_list             (isFC_list_1_3),
    .FCdn_list             (FCdn_list_1_3),
    .FCpl_list             (FCpl_list_1_3),
    .rt_file_list          (cast_rt_file_list_1_3)
)router_1_3(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_30_to_31),
    .west_valid_i          (valid_30_to_31),
    .west_ready_o          (ready_31_to_30),
    .west_data_o           (data_31_to_30),
    .west_valid_o          (valid_31_to_30),
    .west_ready_i          (ready_30_to_31),
    .east_data_i           (data_32_to_31),
    .east_valid_i          (valid_32_to_31),
    .east_ready_o          (ready_31_to_32),
    .east_data_o           (data_31_to_32),
    .east_valid_o          (valid_31_to_32),
    .east_ready_i          (ready_32_to_31),
    .vert0_data_i          (data_21_to_31_v0),
    .vert0_valid_i         (valid_21_to_31_v0),
    .vert0_ready_o         (ready_31_to_21_v0),
    .vert0_data_o          (data_31_to_41_v0),
    .vert0_valid_o         (valid_31_to_41_v0),
    .vert0_ready_i         (ready_41_to_31_v0),
    .vert1_data_i          (data_21_to_31_v1),
    .vert1_valid_i         (valid_21_to_31_v1),
    .vert1_ready_o         (ready_31_to_21_v1),
    .vert1_data_o          (data_31_to_41_v1),
    .vert1_valid_o         (valid_31_to_41_v1),
    .vert1_ready_i         (ready_41_to_31_v1),
    .local_data_i          (data_i[1][3]),
    .local_valid_i         (valid_i[1][3]),
    .local_ready_o         (ready_o[1][3]),
    .local_data_o          (data_o[1][3]),
    .local_valid_o         (valid_o[1][3]),
    .local_ready_i         (ready_i[1][3]),
    .credit_upd            (credit_upd)
);

/*Router 1,4*/    
cast_router #(
    .isUBM_list            (isUBM_list_1_4),
    .isFC_list             (isFC_list_1_4),
    .FCdn_list             (FCdn_list_1_4),
    .FCpl_list             (FCpl_list_1_4),
    .rt_file_list          (cast_rt_file_list_1_4)
)router_1_4(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_40_to_41),
    .west_valid_i          (valid_40_to_41),
    .west_ready_o          (ready_41_to_40),
    .west_data_o           (data_41_to_40),
    .west_valid_o          (valid_41_to_40),
    .west_ready_i          (ready_40_to_41),
    .east_data_i           (data_42_to_41),
    .east_valid_i          (valid_42_to_41),
    .east_ready_o          (ready_41_to_42),
    .east_data_o           (data_41_to_42),
    .east_valid_o          (valid_41_to_42),
    .east_ready_i          (ready_42_to_41),
    .vert0_data_i          (data_31_to_41_v0),
    .vert0_valid_i         (valid_31_to_41_v0),
    .vert0_ready_o         (ready_41_to_31_v0),
    .vert0_data_o          (data_41_to_51_v0),
    .vert0_valid_o         (valid_41_to_51_v0),
    .vert0_ready_i         (ready_51_to_41_v0),
    .vert1_data_i          (data_31_to_41_v1),
    .vert1_valid_i         (valid_31_to_41_v1),
    .vert1_ready_o         (ready_41_to_31_v1),
    .vert1_data_o          (data_41_to_51_v1),
    .vert1_valid_o         (valid_41_to_51_v1),
    .vert1_ready_i         (ready_51_to_41_v1),
    .local_data_i          (data_i[1][4]),
    .local_valid_i         (valid_i[1][4]),
    .local_ready_o         (ready_o[1][4]),
    .local_data_o          (data_o[1][4]),
    .local_valid_o         (valid_o[1][4]),
    .local_ready_i         (ready_i[1][4]),
    .credit_upd            (credit_upd)
);

/*Router 1,5*/    
cast_router #(
    .isUBM_list            (isUBM_list_1_5),
    .isFC_list             (isFC_list_1_5),
    .FCdn_list             (FCdn_list_1_5),
    .FCpl_list             (FCpl_list_1_5),
    .rt_file_list          (cast_rt_file_list_1_5)
)router_1_5(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_50_to_51),
    .west_valid_i          (valid_50_to_51),
    .west_ready_o          (ready_51_to_50),
    .west_data_o           (data_51_to_50),
    .west_valid_o          (valid_51_to_50),
    .west_ready_i          (ready_50_to_51),
    .east_data_i           (data_52_to_51),
    .east_valid_i          (valid_52_to_51),
    .east_ready_o          (ready_51_to_52),
    .east_data_o           (data_51_to_52),
    .east_valid_o          (valid_51_to_52),
    .east_ready_i          (ready_52_to_51),
    .vert0_data_i          (data_41_to_51_v0),
    .vert0_valid_i         (valid_41_to_51_v0),
    .vert0_ready_o         (ready_51_to_41_v0),
    .vert0_data_o          (data_51_to_61_v0),
    .vert0_valid_o         (valid_51_to_61_v0),
    .vert0_ready_i         (ready_61_to_51_v0),
    .vert1_data_i          (data_41_to_51_v1),
    .vert1_valid_i         (valid_41_to_51_v1),
    .vert1_ready_o         (ready_51_to_41_v1),
    .vert1_data_o          (data_51_to_61_v1),
    .vert1_valid_o         (valid_51_to_61_v1),
    .vert1_ready_i         (ready_61_to_51_v1),
    .local_data_i          (data_i[1][5]),
    .local_valid_i         (valid_i[1][5]),
    .local_ready_o         (ready_o[1][5]),
    .local_data_o          (data_o[1][5]),
    .local_valid_o         (valid_o[1][5]),
    .local_ready_i         (ready_i[1][5]),
    .credit_upd            (credit_upd)
);

/*Router 1,6*/    
cast_router #(
    .isUBM_list            (isUBM_list_1_6),
    .isFC_list             (isFC_list_1_6),
    .FCdn_list             (FCdn_list_1_6),
    .FCpl_list             (FCpl_list_1_6),
    .rt_file_list          (cast_rt_file_list_1_6)
)router_1_6(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_60_to_61),
    .west_valid_i          (valid_60_to_61),
    .west_ready_o          (ready_61_to_60),
    .west_data_o           (data_61_to_60),
    .west_valid_o          (valid_61_to_60),
    .west_ready_i          (ready_60_to_61),
    .east_data_i           (data_62_to_61),
    .east_valid_i          (valid_62_to_61),
    .east_ready_o          (ready_61_to_62),
    .east_data_o           (data_61_to_62),
    .east_valid_o          (valid_61_to_62),
    .east_ready_i          (ready_62_to_61),
    .vert0_data_i          (data_51_to_61_v0),
    .vert0_valid_i         (valid_51_to_61_v0),
    .vert0_ready_o         (ready_61_to_51_v0),
    .vert0_data_o          (data_61_to_71_v0),
    .vert0_valid_o         (valid_61_to_71_v0),
    .vert0_ready_i         (ready_71_to_61_v0),
    .vert1_data_i          (data_51_to_61_v1),
    .vert1_valid_i         (valid_51_to_61_v1),
    .vert1_ready_o         (ready_61_to_51_v1),
    .vert1_data_o          (data_61_to_71_v1),
    .vert1_valid_o         (valid_61_to_71_v1),
    .vert1_ready_i         (ready_71_to_61_v1),
    .local_data_i          (data_i[1][6]),
    .local_valid_i         (valid_i[1][6]),
    .local_ready_o         (ready_o[1][6]),
    .local_data_o          (data_o[1][6]),
    .local_valid_o         (valid_o[1][6]),
    .local_ready_i         (ready_i[1][6]),
    .credit_upd            (credit_upd)
);

/*Router 1,7*/    
cast_router #(
    .isUBM_list            (isUBM_list_1_7),
    .isFC_list             (isFC_list_1_7),
    .FCdn_list             (FCdn_list_1_7),
    .FCpl_list             (FCpl_list_1_7),
    .rt_file_list          (cast_rt_file_list_1_7)
)router_1_7(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_70_to_71),
    .west_valid_i          (valid_70_to_71),
    .west_ready_o          (ready_71_to_70),
    .west_data_o           (data_71_to_70),
    .west_valid_o          (valid_71_to_70),
    .west_ready_i          (ready_70_to_71),
    .east_data_i           (data_72_to_71),
    .east_valid_i          (valid_72_to_71),
    .east_ready_o          (ready_71_to_72),
    .east_data_o           (data_71_to_72),
    .east_valid_o          (valid_71_to_72),
    .east_ready_i          (ready_72_to_71),
    .vert0_data_i          (data_61_to_71_v0),
    .vert0_valid_i         (valid_61_to_71_v0),
    .vert0_ready_o         (ready_71_to_61_v0),
    .vert0_data_o          (data_71_to_81_v0),
    .vert0_valid_o         (valid_71_to_81_v0),
    .vert0_ready_i         (ready_81_to_71_v0),
    .vert1_data_i          (data_61_to_71_v1),
    .vert1_valid_i         (valid_61_to_71_v1),
    .vert1_ready_o         (ready_71_to_61_v1),
    .vert1_data_o          (data_71_to_81_v1),
    .vert1_valid_o         (valid_71_to_81_v1),
    .vert1_ready_i         (ready_81_to_71_v1),
    .local_data_i          (data_i[1][7]),
    .local_valid_i         (valid_i[1][7]),
    .local_ready_o         (ready_o[1][7]),
    .local_data_o          (data_o[1][7]),
    .local_valid_o         (valid_o[1][7]),
    .local_ready_i         (ready_i[1][7]),
    .credit_upd            (credit_upd)
);

/*Router 1,8*/    
cast_router #(
    .isUBM_list            (isUBM_list_1_8),
    .isFC_list             (isFC_list_1_8),
    .FCdn_list             (FCdn_list_1_8),
    .FCpl_list             (FCpl_list_1_8),
    .rt_file_list          (cast_rt_file_list_1_8)
)router_1_8(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_80_to_81),
    .west_valid_i          (valid_80_to_81),
    .west_ready_o          (ready_81_to_80),
    .west_data_o           (data_81_to_80),
    .west_valid_o          (valid_81_to_80),
    .west_ready_i          (ready_80_to_81),
    .east_data_i           (data_82_to_81),
    .east_valid_i          (valid_82_to_81),
    .east_ready_o          (ready_81_to_82),
    .east_data_o           (data_81_to_82),
    .east_valid_o          (valid_81_to_82),
    .east_ready_i          (ready_82_to_81),
    .vert0_data_i          (data_71_to_81_v0),
    .vert0_valid_i         (valid_71_to_81_v0),
    .vert0_ready_o         (ready_81_to_71_v0),
    .vert0_data_o          (data_81_to_91_v0),
    .vert0_valid_o         (valid_81_to_91_v0),
    .vert0_ready_i         (ready_91_to_81_v0),
    .vert1_data_i          (data_71_to_81_v1),
    .vert1_valid_i         (valid_71_to_81_v1),
    .vert1_ready_o         (ready_81_to_71_v1),
    .vert1_data_o          (data_81_to_91_v1),
    .vert1_valid_o         (valid_81_to_91_v1),
    .vert1_ready_i         (ready_91_to_81_v1),
    .local_data_i          (data_i[1][8]),
    .local_valid_i         (valid_i[1][8]),
    .local_ready_o         (ready_o[1][8]),
    .local_data_o          (data_o[1][8]),
    .local_valid_o         (valid_o[1][8]),
    .local_ready_i         (ready_i[1][8]),
    .credit_upd            (credit_upd)
);

/*Router 1,9*/    
cast_router #(
    .isUBM_list            (isUBM_list_1_9),
    .isFC_list             (isFC_list_1_9),
    .FCdn_list             (FCdn_list_1_9),
    .FCpl_list             (FCpl_list_1_9),
    .rt_file_list          (cast_rt_file_list_1_9)
)router_1_9(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_90_to_91),
    .west_valid_i          (valid_90_to_91),
    .west_ready_o          (ready_91_to_90),
    .west_data_o           (data_91_to_90),
    .west_valid_o          (valid_91_to_90),
    .west_ready_i          (ready_90_to_91),
    .east_data_i           (data_92_to_91),
    .east_valid_i          (valid_92_to_91),
    .east_ready_o          (ready_91_to_92),
    .east_data_o           (data_91_to_92),
    .east_valid_o          (valid_91_to_92),
    .east_ready_i          (ready_92_to_91),
    .vert0_data_i          (data_81_to_91_v0),
    .vert0_valid_i         (valid_81_to_91_v0),
    .vert0_ready_o         (ready_91_to_81_v0),
    .vert0_data_o          (data_91_to_101_v0),
    .vert0_valid_o         (valid_91_to_101_v0),
    .vert0_ready_i         (ready_101_to_91_v0),
    .vert1_data_i          (data_81_to_91_v1),
    .vert1_valid_i         (valid_81_to_91_v1),
    .vert1_ready_o         (ready_91_to_81_v1),
    .vert1_data_o          (data_91_to_101_v1),
    .vert1_valid_o         (valid_91_to_101_v1),
    .vert1_ready_i         (ready_101_to_91_v1),
    .local_data_i          (data_i[1][9]),
    .local_valid_i         (valid_i[1][9]),
    .local_ready_o         (ready_o[1][9]),
    .local_data_o          (data_o[1][9]),
    .local_valid_o         (valid_o[1][9]),
    .local_ready_i         (ready_i[1][9]),
    .credit_upd            (credit_upd)
);

/*Router 1,10*/    
cast_router #(
    .isUBM_list            (isUBM_list_1_10),
    .isFC_list             (isFC_list_1_10),
    .FCdn_list             (FCdn_list_1_10),
    .FCpl_list             (FCpl_list_1_10),
    .rt_file_list          (cast_rt_file_list_1_10)
)router_1_10(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_100_to_101),
    .west_valid_i          (valid_100_to_101),
    .west_ready_o          (ready_101_to_100),
    .west_data_o           (data_101_to_100),
    .west_valid_o          (valid_101_to_100),
    .west_ready_i          (ready_100_to_101),
    .east_data_i           (data_102_to_101),
    .east_valid_i          (valid_102_to_101),
    .east_ready_o          (ready_101_to_102),
    .east_data_o           (data_101_to_102),
    .east_valid_o          (valid_101_to_102),
    .east_ready_i          (ready_102_to_101),
    .vert0_data_i          (data_91_to_101_v0),
    .vert0_valid_i         (valid_91_to_101_v0),
    .vert0_ready_o         (ready_101_to_91_v0),
    .vert0_data_o          (data_101_to_111_v0),
    .vert0_valid_o         (valid_101_to_111_v0),
    .vert0_ready_i         (ready_111_to_101_v0),
    .vert1_data_i          (data_91_to_101_v1),
    .vert1_valid_i         (valid_91_to_101_v1),
    .vert1_ready_o         (ready_101_to_91_v1),
    .vert1_data_o          (data_101_to_111_v1),
    .vert1_valid_o         (valid_101_to_111_v1),
    .vert1_ready_i         (ready_111_to_101_v1),
    .local_data_i          (data_i[1][10]),
    .local_valid_i         (valid_i[1][10]),
    .local_ready_o         (ready_o[1][10]),
    .local_data_o          (data_o[1][10]),
    .local_valid_o         (valid_o[1][10]),
    .local_ready_i         (ready_i[1][10]),
    .credit_upd            (credit_upd)
);

/*Router 1,11*/    
cast_router #(
    .isUBM_list            (isUBM_list_1_11),
    .isFC_list             (isFC_list_1_11),
    .FCdn_list             (FCdn_list_1_11),
    .FCpl_list             (FCpl_list_1_11),
    .rt_file_list          (cast_rt_file_list_1_11)
)router_1_11(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_110_to_111),
    .west_valid_i          (valid_110_to_111),
    .west_ready_o          (ready_111_to_110),
    .west_data_o           (data_111_to_110),
    .west_valid_o          (valid_111_to_110),
    .west_ready_i          (ready_110_to_111),
    .east_data_i           (data_112_to_111),
    .east_valid_i          (valid_112_to_111),
    .east_ready_o          (ready_111_to_112),
    .east_data_o           (data_111_to_112),
    .east_valid_o          (valid_111_to_112),
    .east_ready_i          (ready_112_to_111),
    .vert0_data_i          (data_101_to_111_v0),
    .vert0_valid_i         (valid_101_to_111_v0),
    .vert0_ready_o         (ready_111_to_101_v0),
    .vert0_data_o          (data_111_to_121_v0),
    .vert0_valid_o         (valid_111_to_121_v0),
    .vert0_ready_i         (ready_121_to_111_v0),
    .vert1_data_i          (data_101_to_111_v1),
    .vert1_valid_i         (valid_101_to_111_v1),
    .vert1_ready_o         (ready_111_to_101_v1),
    .vert1_data_o          (data_111_to_121_v1),
    .vert1_valid_o         (valid_111_to_121_v1),
    .vert1_ready_i         (ready_121_to_111_v1),
    .local_data_i          (data_i[1][11]),
    .local_valid_i         (valid_i[1][11]),
    .local_ready_o         (ready_o[1][11]),
    .local_data_o          (data_o[1][11]),
    .local_valid_o         (valid_o[1][11]),
    .local_ready_i         (ready_i[1][11]),
    .credit_upd            (credit_upd)
);

/*Router 1,12*/    
cast_router #(
    .isUBM_list            (isUBM_list_1_12),
    .isFC_list             (isFC_list_1_12),
    .FCdn_list             (FCdn_list_1_12),
    .FCpl_list             (FCpl_list_1_12),
    .rt_file_list          (cast_rt_file_list_1_12)
)router_1_12(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_120_to_121),
    .west_valid_i          (valid_120_to_121),
    .west_ready_o          (ready_121_to_120),
    .west_data_o           (data_121_to_120),
    .west_valid_o          (valid_121_to_120),
    .west_ready_i          (ready_120_to_121),
    .east_data_i           (data_122_to_121),
    .east_valid_i          (valid_122_to_121),
    .east_ready_o          (ready_121_to_122),
    .east_data_o           (data_121_to_122),
    .east_valid_o          (valid_121_to_122),
    .east_ready_i          (ready_122_to_121),
    .vert0_data_i          (data_111_to_121_v0),
    .vert0_valid_i         (valid_111_to_121_v0),
    .vert0_ready_o         (ready_121_to_111_v0),
    .vert0_data_o          (data_121_to_131_v0),
    .vert0_valid_o         (valid_121_to_131_v0),
    .vert0_ready_i         (ready_131_to_121_v0),
    .vert1_data_i          (data_111_to_121_v1),
    .vert1_valid_i         (valid_111_to_121_v1),
    .vert1_ready_o         (ready_121_to_111_v1),
    .vert1_data_o          (data_121_to_131_v1),
    .vert1_valid_o         (valid_121_to_131_v1),
    .vert1_ready_i         (ready_131_to_121_v1),
    .local_data_i          (data_i[1][12]),
    .local_valid_i         (valid_i[1][12]),
    .local_ready_o         (ready_o[1][12]),
    .local_data_o          (data_o[1][12]),
    .local_valid_o         (valid_o[1][12]),
    .local_ready_i         (ready_i[1][12]),
    .credit_upd            (credit_upd)
);

/*Router 1,13*/    
cast_router #(
    .isUBM_list            (isUBM_list_1_13),
    .isFC_list             (isFC_list_1_13),
    .FCdn_list             (FCdn_list_1_13),
    .FCpl_list             (FCpl_list_1_13),
    .rt_file_list          (cast_rt_file_list_1_13)
)router_1_13(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_130_to_131),
    .west_valid_i          (valid_130_to_131),
    .west_ready_o          (ready_131_to_130),
    .west_data_o           (data_131_to_130),
    .west_valid_o          (valid_131_to_130),
    .west_ready_i          (ready_130_to_131),
    .east_data_i           (data_132_to_131),
    .east_valid_i          (valid_132_to_131),
    .east_ready_o          (ready_131_to_132),
    .east_data_o           (data_131_to_132),
    .east_valid_o          (valid_131_to_132),
    .east_ready_i          (ready_132_to_131),
    .vert0_data_i          (data_121_to_131_v0),
    .vert0_valid_i         (valid_121_to_131_v0),
    .vert0_ready_o         (ready_131_to_121_v0),
    .vert0_data_o          (data_131_to_141_v0),
    .vert0_valid_o         (valid_131_to_141_v0),
    .vert0_ready_i         (ready_141_to_131_v0),
    .vert1_data_i          (data_121_to_131_v1),
    .vert1_valid_i         (valid_121_to_131_v1),
    .vert1_ready_o         (ready_131_to_121_v1),
    .vert1_data_o          (data_131_to_141_v1),
    .vert1_valid_o         (valid_131_to_141_v1),
    .vert1_ready_i         (ready_141_to_131_v1),
    .local_data_i          (data_i[1][13]),
    .local_valid_i         (valid_i[1][13]),
    .local_ready_o         (ready_o[1][13]),
    .local_data_o          (data_o[1][13]),
    .local_valid_o         (valid_o[1][13]),
    .local_ready_i         (ready_i[1][13]),
    .credit_upd            (credit_upd)
);

/*Router 1,14*/    
cast_router #(
    .isUBM_list            (isUBM_list_1_14),
    .isFC_list             (isFC_list_1_14),
    .FCdn_list             (FCdn_list_1_14),
    .FCpl_list             (FCpl_list_1_14),
    .rt_file_list          (cast_rt_file_list_1_14)
)router_1_14(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_140_to_141),
    .west_valid_i          (valid_140_to_141),
    .west_ready_o          (ready_141_to_140),
    .west_data_o           (data_141_to_140),
    .west_valid_o          (valid_141_to_140),
    .west_ready_i          (ready_140_to_141),
    .east_data_i           (data_142_to_141),
    .east_valid_i          (valid_142_to_141),
    .east_ready_o          (ready_141_to_142),
    .east_data_o           (data_141_to_142),
    .east_valid_o          (valid_141_to_142),
    .east_ready_i          (ready_142_to_141),
    .vert0_data_i          (data_131_to_141_v0),
    .vert0_valid_i         (valid_131_to_141_v0),
    .vert0_ready_o         (ready_141_to_131_v0),
    .vert0_data_o          (data_141_to_151_v0),
    .vert0_valid_o         (valid_141_to_151_v0),
    .vert0_ready_i         (ready_151_to_141_v0),
    .vert1_data_i          (data_131_to_141_v1),
    .vert1_valid_i         (valid_131_to_141_v1),
    .vert1_ready_o         (ready_141_to_131_v1),
    .vert1_data_o          (data_141_to_151_v1),
    .vert1_valid_o         (valid_141_to_151_v1),
    .vert1_ready_i         (ready_151_to_141_v1),
    .local_data_i          (data_i[1][14]),
    .local_valid_i         (valid_i[1][14]),
    .local_ready_o         (ready_o[1][14]),
    .local_data_o          (data_o[1][14]),
    .local_valid_o         (valid_o[1][14]),
    .local_ready_i         (ready_i[1][14]),
    .credit_upd            (credit_upd)
);

/*Router 1,15*/    
cast_router #(
    .isUBM_list            (isUBM_list_1_15),
    .isFC_list             (isFC_list_1_15),
    .FCdn_list             (FCdn_list_1_15),
    .FCpl_list             (FCpl_list_1_15),
    .rt_file_list          (cast_rt_file_list_1_15)
)router_1_15(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_150_to_151),
    .west_valid_i          (valid_150_to_151),
    .west_ready_o          (ready_151_to_150),
    .west_data_o           (data_151_to_150),
    .west_valid_o          (valid_151_to_150),
    .west_ready_i          (ready_150_to_151),
    .east_data_i           (data_152_to_151),
    .east_valid_i          (valid_152_to_151),
    .east_ready_o          (ready_151_to_152),
    .east_data_o           (data_151_to_152),
    .east_valid_o          (valid_151_to_152),
    .east_ready_i          (ready_152_to_151),
    .vert0_data_i          (data_141_to_151_v0),
    .vert0_valid_i         (valid_141_to_151_v0),
    .vert0_ready_o         (ready_151_to_141_v0),
    .vert0_data_o          (data_151_to_161_v0),
    .vert0_valid_o         (valid_151_to_161_v0),
    .vert0_ready_i         (ready_161_to_151_v0),
    .vert1_data_i          (data_141_to_151_v1),
    .vert1_valid_i         (valid_141_to_151_v1),
    .vert1_ready_o         (ready_151_to_141_v1),
    .vert1_data_o          (data_151_to_161_v1),
    .vert1_valid_o         (valid_151_to_161_v1),
    .vert1_ready_i         (ready_161_to_151_v1),
    .local_data_i          (data_i[1][15]),
    .local_valid_i         (valid_i[1][15]),
    .local_ready_o         (ready_o[1][15]),
    .local_data_o          (data_o[1][15]),
    .local_valid_o         (valid_o[1][15]),
    .local_ready_i         (ready_i[1][15]),
    .credit_upd            (credit_upd)
);

/*Router 1,16*/    
cast_router #(
    .isUBM_list            (isUBM_list_1_16),
    .isFC_list             (isFC_list_1_16),
    .FCdn_list             (FCdn_list_1_16),
    .FCpl_list             (FCpl_list_1_16),
    .rt_file_list          (cast_rt_file_list_1_16)
)router_1_16(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_160_to_161),
    .west_valid_i          (valid_160_to_161),
    .west_ready_o          (ready_161_to_160),
    .west_data_o           (data_161_to_160),
    .west_valid_o          (valid_161_to_160),
    .west_ready_i          (ready_160_to_161),
    .east_data_i           (data_162_to_161),
    .east_valid_i          (valid_162_to_161),
    .east_ready_o          (ready_161_to_162),
    .east_data_o           (data_161_to_162),
    .east_valid_o          (valid_161_to_162),
    .east_ready_i          (ready_162_to_161),
    .vert0_data_i          (data_151_to_161_v0),
    .vert0_valid_i         (valid_151_to_161_v0),
    .vert0_ready_o         (ready_161_to_151_v0),
    .vert0_data_o          (data_161_to_171_v0),
    .vert0_valid_o         (valid_161_to_171_v0),
    .vert0_ready_i         (ready_171_to_161_v0),
    .vert1_data_i          (data_151_to_161_v1),
    .vert1_valid_i         (valid_151_to_161_v1),
    .vert1_ready_o         (ready_161_to_151_v1),
    .vert1_data_o          (data_161_to_171_v1),
    .vert1_valid_o         (valid_161_to_171_v1),
    .vert1_ready_i         (ready_171_to_161_v1),
    .local_data_i          (data_i[1][16]),
    .local_valid_i         (valid_i[1][16]),
    .local_ready_o         (ready_o[1][16]),
    .local_data_o          (data_o[1][16]),
    .local_valid_o         (valid_o[1][16]),
    .local_ready_i         (ready_i[1][16]),
    .credit_upd            (credit_upd)
);

/*Router 1,17*/    
cast_router #(
    .isUBM_list            (isUBM_list_1_17),
    .isFC_list             (isFC_list_1_17),
    .FCdn_list             (FCdn_list_1_17),
    .FCpl_list             (FCpl_list_1_17),
    .rt_file_list          (cast_rt_file_list_1_17)
)router_1_17(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_170_to_171),
    .west_valid_i          (valid_170_to_171),
    .west_ready_o          (ready_171_to_170),
    .west_data_o           (data_171_to_170),
    .west_valid_o          (valid_171_to_170),
    .west_ready_i          (ready_170_to_171),
    .east_data_i           (data_172_to_171),
    .east_valid_i          (valid_172_to_171),
    .east_ready_o          (ready_171_to_172),
    .east_data_o           (data_171_to_172),
    .east_valid_o          (valid_171_to_172),
    .east_ready_i          (ready_172_to_171),
    .vert0_data_i          (data_161_to_171_v0),
    .vert0_valid_i         (valid_161_to_171_v0),
    .vert0_ready_o         (ready_171_to_161_v0),
    .vert0_data_o          (data_171_to_181_v0),
    .vert0_valid_o         (valid_171_to_181_v0),
    .vert0_ready_i         (ready_181_to_171_v0),
    .vert1_data_i          (data_161_to_171_v1),
    .vert1_valid_i         (valid_161_to_171_v1),
    .vert1_ready_o         (ready_171_to_161_v1),
    .vert1_data_o          (data_171_to_181_v1),
    .vert1_valid_o         (valid_171_to_181_v1),
    .vert1_ready_i         (ready_181_to_171_v1),
    .local_data_i          (data_i[1][17]),
    .local_valid_i         (valid_i[1][17]),
    .local_ready_o         (ready_o[1][17]),
    .local_data_o          (data_o[1][17]),
    .local_valid_o         (valid_o[1][17]),
    .local_ready_i         (ready_i[1][17]),
    .credit_upd            (credit_upd)
);

/*Router 1,18*/    
cast_router #(
    .isUBM_list            (isUBM_list_1_18),
    .isFC_list             (isFC_list_1_18),
    .FCdn_list             (FCdn_list_1_18),
    .FCpl_list             (FCpl_list_1_18),
    .rt_file_list          (cast_rt_file_list_1_18)
)router_1_18(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_180_to_181),
    .west_valid_i          (valid_180_to_181),
    .west_ready_o          (ready_181_to_180),
    .west_data_o           (data_181_to_180),
    .west_valid_o          (valid_181_to_180),
    .west_ready_i          (ready_180_to_181),
    .east_data_i           (data_182_to_181),
    .east_valid_i          (valid_182_to_181),
    .east_ready_o          (ready_181_to_182),
    .east_data_o           (data_181_to_182),
    .east_valid_o          (valid_181_to_182),
    .east_ready_i          (ready_182_to_181),
    .vert0_data_i          (data_171_to_181_v0),
    .vert0_valid_i         (valid_171_to_181_v0),
    .vert0_ready_o         (ready_181_to_171_v0),
    .vert0_data_o          (data_181_to_191_v0),
    .vert0_valid_o         (valid_181_to_191_v0),
    .vert0_ready_i         (ready_191_to_181_v0),
    .vert1_data_i          (data_171_to_181_v1),
    .vert1_valid_i         (valid_171_to_181_v1),
    .vert1_ready_o         (ready_181_to_171_v1),
    .vert1_data_o          (data_181_to_191_v1),
    .vert1_valid_o         (valid_181_to_191_v1),
    .vert1_ready_i         (ready_191_to_181_v1),
    .local_data_i          (data_i[1][18]),
    .local_valid_i         (valid_i[1][18]),
    .local_ready_o         (ready_o[1][18]),
    .local_data_o          (data_o[1][18]),
    .local_valid_o         (valid_o[1][18]),
    .local_ready_i         (ready_i[1][18]),
    .credit_upd            (credit_upd)
);

/*Router 1,19*/    
cast_router #(
    .isUBM_list            (isUBM_list_1_19),
    .isFC_list             (isFC_list_1_19),
    .FCdn_list             (FCdn_list_1_19),
    .FCpl_list             (FCpl_list_1_19),
    .rt_file_list          (cast_rt_file_list_1_19)
)router_1_19(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_190_to_191),
    .west_valid_i          (valid_190_to_191),
    .west_ready_o          (ready_191_to_190),
    .west_data_o           (data_191_to_190),
    .west_valid_o          (valid_191_to_190),
    .west_ready_i          (ready_190_to_191),
    .east_data_i           (data_192_to_191),
    .east_valid_i          (valid_192_to_191),
    .east_ready_o          (ready_191_to_192),
    .east_data_o           (data_191_to_192),
    .east_valid_o          (valid_191_to_192),
    .east_ready_i          (ready_192_to_191),
    .vert0_data_i          (data_181_to_191_v0),
    .vert0_valid_i         (valid_181_to_191_v0),
    .vert0_ready_o         (ready_191_to_181_v0),
    .vert0_data_o          (data_191_to_201_v0),
    .vert0_valid_o         (valid_191_to_201_v0),
    .vert0_ready_i         (ready_201_to_191_v0),
    .vert1_data_i          (data_181_to_191_v1),
    .vert1_valid_i         (valid_181_to_191_v1),
    .vert1_ready_o         (ready_191_to_181_v1),
    .vert1_data_o          (data_191_to_201_v1),
    .vert1_valid_o         (valid_191_to_201_v1),
    .vert1_ready_i         (ready_201_to_191_v1),
    .local_data_i          (data_i[1][19]),
    .local_valid_i         (valid_i[1][19]),
    .local_ready_o         (ready_o[1][19]),
    .local_data_o          (data_o[1][19]),
    .local_valid_o         (valid_o[1][19]),
    .local_ready_i         (ready_i[1][19]),
    .credit_upd            (credit_upd)
);

/*Router 1,20*/    
cast_router #(
    .isUBM_list            (isUBM_list_1_20),
    .isFC_list             (isFC_list_1_20),
    .FCdn_list             (FCdn_list_1_20),
    .FCpl_list             (FCpl_list_1_20),
    .rt_file_list          (cast_rt_file_list_1_20)
)router_1_20(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_200_to_201),
    .west_valid_i          (valid_200_to_201),
    .west_ready_o          (ready_201_to_200),
    .west_data_o           (data_201_to_200),
    .west_valid_o          (valid_201_to_200),
    .west_ready_i          (ready_200_to_201),
    .east_data_i           (data_202_to_201),
    .east_valid_i          (valid_202_to_201),
    .east_ready_o          (ready_201_to_202),
    .east_data_o           (data_201_to_202),
    .east_valid_o          (valid_201_to_202),
    .east_ready_i          (ready_202_to_201),
    .vert0_data_i          (data_191_to_201_v0),
    .vert0_valid_i         (valid_191_to_201_v0),
    .vert0_ready_o         (ready_201_to_191_v0),
    .vert0_data_o          (data_201_to_211_v0),
    .vert0_valid_o         (valid_201_to_211_v0),
    .vert0_ready_i         (ready_211_to_201_v0),
    .vert1_data_i          (data_191_to_201_v1),
    .vert1_valid_i         (valid_191_to_201_v1),
    .vert1_ready_o         (ready_201_to_191_v1),
    .vert1_data_o          (data_201_to_211_v1),
    .vert1_valid_o         (valid_201_to_211_v1),
    .vert1_ready_i         (ready_211_to_201_v1),
    .local_data_i          (data_i[1][20]),
    .local_valid_i         (valid_i[1][20]),
    .local_ready_o         (ready_o[1][20]),
    .local_data_o          (data_o[1][20]),
    .local_valid_o         (valid_o[1][20]),
    .local_ready_i         (ready_i[1][20]),
    .credit_upd            (credit_upd)
);

/*Router 1,21*/    
cast_router #(
    .isUBM_list            (isUBM_list_1_21),
    .isFC_list             (isFC_list_1_21),
    .FCdn_list             (FCdn_list_1_21),
    .FCpl_list             (FCpl_list_1_21),
    .rt_file_list          (cast_rt_file_list_1_21)
)router_1_21(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_210_to_211),
    .west_valid_i          (valid_210_to_211),
    .west_ready_o          (ready_211_to_210),
    .west_data_o           (data_211_to_210),
    .west_valid_o          (valid_211_to_210),
    .west_ready_i          (ready_210_to_211),
    .east_data_i           (data_212_to_211),
    .east_valid_i          (valid_212_to_211),
    .east_ready_o          (ready_211_to_212),
    .east_data_o           (data_211_to_212),
    .east_valid_o          (valid_211_to_212),
    .east_ready_i          (ready_212_to_211),
    .vert0_data_i          (data_201_to_211_v0),
    .vert0_valid_i         (valid_201_to_211_v0),
    .vert0_ready_o         (ready_211_to_201_v0),
    .vert0_data_o          (data_211_to_221_v0),
    .vert0_valid_o         (valid_211_to_221_v0),
    .vert0_ready_i         (ready_221_to_211_v0),
    .vert1_data_i          (data_201_to_211_v1),
    .vert1_valid_i         (valid_201_to_211_v1),
    .vert1_ready_o         (ready_211_to_201_v1),
    .vert1_data_o          (data_211_to_221_v1),
    .vert1_valid_o         (valid_211_to_221_v1),
    .vert1_ready_i         (ready_221_to_211_v1),
    .local_data_i          (data_i[1][21]),
    .local_valid_i         (valid_i[1][21]),
    .local_ready_o         (ready_o[1][21]),
    .local_data_o          (data_o[1][21]),
    .local_valid_o         (valid_o[1][21]),
    .local_ready_i         (ready_i[1][21]),
    .credit_upd            (credit_upd)
);

/*Router 1,22*/    
cast_router #(
    .isUBM_list            (isUBM_list_1_22),
    .isFC_list             (isFC_list_1_22),
    .FCdn_list             (FCdn_list_1_22),
    .FCpl_list             (FCpl_list_1_22),
    .rt_file_list          (cast_rt_file_list_1_22)
)router_1_22(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_220_to_221),
    .west_valid_i          (valid_220_to_221),
    .west_ready_o          (ready_221_to_220),
    .west_data_o           (data_221_to_220),
    .west_valid_o          (valid_221_to_220),
    .west_ready_i          (ready_220_to_221),
    .east_data_i           (data_222_to_221),
    .east_valid_i          (valid_222_to_221),
    .east_ready_o          (ready_221_to_222),
    .east_data_o           (data_221_to_222),
    .east_valid_o          (valid_221_to_222),
    .east_ready_i          (ready_222_to_221),
    .vert0_data_i          (data_211_to_221_v0),
    .vert0_valid_i         (valid_211_to_221_v0),
    .vert0_ready_o         (ready_221_to_211_v0),
    .vert0_data_o          (data_221_to_231_v0),
    .vert0_valid_o         (valid_221_to_231_v0),
    .vert0_ready_i         (ready_231_to_221_v0),
    .vert1_data_i          (data_211_to_221_v1),
    .vert1_valid_i         (valid_211_to_221_v1),
    .vert1_ready_o         (ready_221_to_211_v1),
    .vert1_data_o          (data_221_to_231_v1),
    .vert1_valid_o         (valid_221_to_231_v1),
    .vert1_ready_i         (ready_231_to_221_v1),
    .local_data_i          (data_i[1][22]),
    .local_valid_i         (valid_i[1][22]),
    .local_ready_o         (ready_o[1][22]),
    .local_data_o          (data_o[1][22]),
    .local_valid_o         (valid_o[1][22]),
    .local_ready_i         (ready_i[1][22]),
    .credit_upd            (credit_upd)
);

/*Router 1,23*/    
cast_router #(
    .isUBM_list            (isUBM_list_1_23),
    .isFC_list             (isFC_list_1_23),
    .FCdn_list             (FCdn_list_1_23),
    .FCpl_list             (FCpl_list_1_23),
    .rt_file_list          (cast_rt_file_list_1_23)
)router_1_23(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_230_to_231),
    .west_valid_i          (valid_230_to_231),
    .west_ready_o          (ready_231_to_230),
    .west_data_o           (data_231_to_230),
    .west_valid_o          (valid_231_to_230),
    .west_ready_i          (ready_230_to_231),
    .east_data_i           (data_232_to_231),
    .east_valid_i          (valid_232_to_231),
    .east_ready_o          (ready_231_to_232),
    .east_data_o           (data_231_to_232),
    .east_valid_o          (valid_231_to_232),
    .east_ready_i          (ready_232_to_231),
    .vert0_data_i          (data_221_to_231_v0),
    .vert0_valid_i         (valid_221_to_231_v0),
    .vert0_ready_o         (ready_231_to_221_v0),
    .vert0_data_o          (data_231_to_241_v0),
    .vert0_valid_o         (valid_231_to_241_v0),
    .vert0_ready_i         (ready_241_to_231_v0),
    .vert1_data_i          (data_221_to_231_v1),
    .vert1_valid_i         (valid_221_to_231_v1),
    .vert1_ready_o         (ready_231_to_221_v1),
    .vert1_data_o          (data_231_to_241_v1),
    .vert1_valid_o         (valid_231_to_241_v1),
    .vert1_ready_i         (ready_241_to_231_v1),
    .local_data_i          (data_i[1][23]),
    .local_valid_i         (valid_i[1][23]),
    .local_ready_o         (ready_o[1][23]),
    .local_data_o          (data_o[1][23]),
    .local_valid_o         (valid_o[1][23]),
    .local_ready_i         (ready_i[1][23]),
    .credit_upd            (credit_upd)
);

/*Router 1,24*/    
cast_router #(
    .isUBM_list            (isUBM_list_1_24),
    .isFC_list             (isFC_list_1_24),
    .FCdn_list             (FCdn_list_1_24),
    .FCpl_list             (FCpl_list_1_24),
    .rt_file_list          (cast_rt_file_list_1_24)
)router_1_24(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_240_to_241),
    .west_valid_i          (valid_240_to_241),
    .west_ready_o          (ready_241_to_240),
    .west_data_o           (data_241_to_240),
    .west_valid_o          (valid_241_to_240),
    .west_ready_i          (ready_240_to_241),
    .east_data_i           (data_242_to_241),
    .east_valid_i          (valid_242_to_241),
    .east_ready_o          (ready_241_to_242),
    .east_data_o           (data_o_flee7),
    .east_valid_o          (valid_o_flee7),
    .east_ready_i          (ready_i_flee7),
    .vert0_data_i          (data_231_to_241_v0),
    .vert0_valid_i         (valid_231_to_241_v0),
    .vert0_ready_o         (ready_241_to_231_v0),
    .vert0_data_o          (),
    .vert0_valid_o         (),
    .vert0_ready_i         (1'b0),
    .vert1_data_i          (data_231_to_241_v1),
    .vert1_valid_i         (valid_231_to_241_v1),
    .vert1_ready_o         (ready_241_to_231_v1),
    .vert1_data_o          (),
    .vert1_valid_o         (),
    .vert1_ready_i         (1'b0),
    .local_data_i          (data_i[1][24]),
    .local_valid_i         (valid_i[1][24]),
    .local_ready_o         (ready_o[1][24]),
    .local_data_o          (data_o[1][24]),
    .local_valid_o         (valid_o[1][24]),
    .local_ready_i         (ready_i[1][24]),
    .credit_upd            (credit_upd)
);

/*Router 2,0*/    
cast_router #(
    .isUBM_list            (isUBM_list_2_0),
    .isFC_list             (isFC_list_2_0),
    .FCdn_list             (FCdn_list_2_0),
    .FCpl_list             (FCpl_list_2_0),
    .rt_file_list          (cast_rt_file_list_2_0)
)router_2_0(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_1_to_2),
    .west_valid_i          (valid_1_to_2),
    .west_ready_o          (ready_2_to_1),
    .west_data_o           (data_2_to_1),
    .west_valid_o          (valid_2_to_1),
    .west_ready_i          (ready_1_to_2),
    .east_data_i           (data_3_to_2),
    .east_valid_i          (valid_3_to_2),
    .east_ready_o          (ready_2_to_3),
    .east_data_o           (data_2_to_3),
    .east_valid_o          (valid_2_to_3),
    .east_ready_i          (ready_3_to_2),
    .vert0_data_i          (34'b0),
    .vert0_valid_i         (1'b0),
    .vert0_ready_o         (),
    .vert0_data_o          (data_2_to_12_v0),
    .vert0_valid_o         (valid_2_to_12_v0),
    .vert0_ready_i         (ready_12_to_2_v0),
    .vert1_data_i          (34'b0),
    .vert1_valid_i         (1'b0),
    .vert1_ready_o         (),
    .vert1_data_o          (data_2_to_12_v1),
    .vert1_valid_o         (valid_2_to_12_v1),
    .vert1_ready_i         (ready_12_to_2_v1),
    .local_data_i          (data_i[2][0]),
    .local_valid_i         (valid_i[2][0]),
    .local_ready_o         (ready_o[2][0]),
    .local_data_o          (data_o[2][0]),
    .local_valid_o         (valid_o[2][0]),
    .local_ready_i         (ready_i[2][0]),
    .credit_upd            (credit_upd)
);

/*Router 2,1*/    
cast_router #(
    .isUBM_list            (isUBM_list_2_1),
    .isFC_list             (isFC_list_2_1),
    .FCdn_list             (FCdn_list_2_1),
    .FCpl_list             (FCpl_list_2_1),
    .rt_file_list          (cast_rt_file_list_2_1)
)router_2_1(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_11_to_12),
    .west_valid_i          (valid_11_to_12),
    .west_ready_o          (ready_12_to_11),
    .west_data_o           (data_12_to_11),
    .west_valid_o          (valid_12_to_11),
    .west_ready_i          (ready_11_to_12),
    .east_data_i           (data_13_to_12),
    .east_valid_i          (valid_13_to_12),
    .east_ready_o          (ready_12_to_13),
    .east_data_o           (data_12_to_13),
    .east_valid_o          (valid_12_to_13),
    .east_ready_i          (ready_13_to_12),
    .vert0_data_i          (data_2_to_12_v0),
    .vert0_valid_i         (valid_2_to_12_v0),
    .vert0_ready_o         (ready_12_to_2_v0),
    .vert0_data_o          (data_12_to_22_v0),
    .vert0_valid_o         (valid_12_to_22_v0),
    .vert0_ready_i         (ready_22_to_12_v0),
    .vert1_data_i          (data_2_to_12_v1),
    .vert1_valid_i         (valid_2_to_12_v1),
    .vert1_ready_o         (ready_12_to_2_v1),
    .vert1_data_o          (data_12_to_22_v1),
    .vert1_valid_o         (valid_12_to_22_v1),
    .vert1_ready_i         (ready_22_to_12_v1),
    .local_data_i          (data_i[2][1]),
    .local_valid_i         (valid_i[2][1]),
    .local_ready_o         (ready_o[2][1]),
    .local_data_o          (data_o[2][1]),
    .local_valid_o         (valid_o[2][1]),
    .local_ready_i         (ready_i[2][1]),
    .credit_upd            (credit_upd)
);

/*Router 2,2*/    
cast_router #(
    .isUBM_list            (isUBM_list_2_2),
    .isFC_list             (isFC_list_2_2),
    .FCdn_list             (FCdn_list_2_2),
    .FCpl_list             (FCpl_list_2_2),
    .rt_file_list          (cast_rt_file_list_2_2)
)router_2_2(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_21_to_22),
    .west_valid_i          (valid_21_to_22),
    .west_ready_o          (ready_22_to_21),
    .west_data_o           (data_22_to_21),
    .west_valid_o          (valid_22_to_21),
    .west_ready_i          (ready_21_to_22),
    .east_data_i           (data_23_to_22),
    .east_valid_i          (valid_23_to_22),
    .east_ready_o          (ready_22_to_23),
    .east_data_o           (data_22_to_23),
    .east_valid_o          (valid_22_to_23),
    .east_ready_i          (ready_23_to_22),
    .vert0_data_i          (data_12_to_22_v0),
    .vert0_valid_i         (valid_12_to_22_v0),
    .vert0_ready_o         (ready_22_to_12_v0),
    .vert0_data_o          (data_22_to_32_v0),
    .vert0_valid_o         (valid_22_to_32_v0),
    .vert0_ready_i         (ready_32_to_22_v0),
    .vert1_data_i          (data_12_to_22_v1),
    .vert1_valid_i         (valid_12_to_22_v1),
    .vert1_ready_o         (ready_22_to_12_v1),
    .vert1_data_o          (data_22_to_32_v1),
    .vert1_valid_o         (valid_22_to_32_v1),
    .vert1_ready_i         (ready_32_to_22_v1),
    .local_data_i          (data_i[2][2]),
    .local_valid_i         (valid_i[2][2]),
    .local_ready_o         (ready_o[2][2]),
    .local_data_o          (data_o[2][2]),
    .local_valid_o         (valid_o[2][2]),
    .local_ready_i         (ready_i[2][2]),
    .credit_upd            (credit_upd)
);

/*Router 2,3*/    
cast_router #(
    .isUBM_list            (isUBM_list_2_3),
    .isFC_list             (isFC_list_2_3),
    .FCdn_list             (FCdn_list_2_3),
    .FCpl_list             (FCpl_list_2_3),
    .rt_file_list          (cast_rt_file_list_2_3)
)router_2_3(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_31_to_32),
    .west_valid_i          (valid_31_to_32),
    .west_ready_o          (ready_32_to_31),
    .west_data_o           (data_32_to_31),
    .west_valid_o          (valid_32_to_31),
    .west_ready_i          (ready_31_to_32),
    .east_data_i           (data_33_to_32),
    .east_valid_i          (valid_33_to_32),
    .east_ready_o          (ready_32_to_33),
    .east_data_o           (data_32_to_33),
    .east_valid_o          (valid_32_to_33),
    .east_ready_i          (ready_33_to_32),
    .vert0_data_i          (data_22_to_32_v0),
    .vert0_valid_i         (valid_22_to_32_v0),
    .vert0_ready_o         (ready_32_to_22_v0),
    .vert0_data_o          (data_32_to_42_v0),
    .vert0_valid_o         (valid_32_to_42_v0),
    .vert0_ready_i         (ready_42_to_32_v0),
    .vert1_data_i          (data_22_to_32_v1),
    .vert1_valid_i         (valid_22_to_32_v1),
    .vert1_ready_o         (ready_32_to_22_v1),
    .vert1_data_o          (data_32_to_42_v1),
    .vert1_valid_o         (valid_32_to_42_v1),
    .vert1_ready_i         (ready_42_to_32_v1),
    .local_data_i          (data_i[2][3]),
    .local_valid_i         (valid_i[2][3]),
    .local_ready_o         (ready_o[2][3]),
    .local_data_o          (data_o[2][3]),
    .local_valid_o         (valid_o[2][3]),
    .local_ready_i         (ready_i[2][3]),
    .credit_upd            (credit_upd)
);

/*Router 2,4*/    
cast_router #(
    .isUBM_list            (isUBM_list_2_4),
    .isFC_list             (isFC_list_2_4),
    .FCdn_list             (FCdn_list_2_4),
    .FCpl_list             (FCpl_list_2_4),
    .rt_file_list          (cast_rt_file_list_2_4)
)router_2_4(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_41_to_42),
    .west_valid_i          (valid_41_to_42),
    .west_ready_o          (ready_42_to_41),
    .west_data_o           (data_42_to_41),
    .west_valid_o          (valid_42_to_41),
    .west_ready_i          (ready_41_to_42),
    .east_data_i           (data_43_to_42),
    .east_valid_i          (valid_43_to_42),
    .east_ready_o          (ready_42_to_43),
    .east_data_o           (data_42_to_43),
    .east_valid_o          (valid_42_to_43),
    .east_ready_i          (ready_43_to_42),
    .vert0_data_i          (data_32_to_42_v0),
    .vert0_valid_i         (valid_32_to_42_v0),
    .vert0_ready_o         (ready_42_to_32_v0),
    .vert0_data_o          (data_42_to_52_v0),
    .vert0_valid_o         (valid_42_to_52_v0),
    .vert0_ready_i         (ready_52_to_42_v0),
    .vert1_data_i          (data_32_to_42_v1),
    .vert1_valid_i         (valid_32_to_42_v1),
    .vert1_ready_o         (ready_42_to_32_v1),
    .vert1_data_o          (data_42_to_52_v1),
    .vert1_valid_o         (valid_42_to_52_v1),
    .vert1_ready_i         (ready_52_to_42_v1),
    .local_data_i          (data_i[2][4]),
    .local_valid_i         (valid_i[2][4]),
    .local_ready_o         (ready_o[2][4]),
    .local_data_o          (data_o[2][4]),
    .local_valid_o         (valid_o[2][4]),
    .local_ready_i         (ready_i[2][4]),
    .credit_upd            (credit_upd)
);

/*Router 2,5*/    
cast_router #(
    .isUBM_list            (isUBM_list_2_5),
    .isFC_list             (isFC_list_2_5),
    .FCdn_list             (FCdn_list_2_5),
    .FCpl_list             (FCpl_list_2_5),
    .rt_file_list          (cast_rt_file_list_2_5)
)router_2_5(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_51_to_52),
    .west_valid_i          (valid_51_to_52),
    .west_ready_o          (ready_52_to_51),
    .west_data_o           (data_52_to_51),
    .west_valid_o          (valid_52_to_51),
    .west_ready_i          (ready_51_to_52),
    .east_data_i           (data_53_to_52),
    .east_valid_i          (valid_53_to_52),
    .east_ready_o          (ready_52_to_53),
    .east_data_o           (data_52_to_53),
    .east_valid_o          (valid_52_to_53),
    .east_ready_i          (ready_53_to_52),
    .vert0_data_i          (data_42_to_52_v0),
    .vert0_valid_i         (valid_42_to_52_v0),
    .vert0_ready_o         (ready_52_to_42_v0),
    .vert0_data_o          (data_52_to_62_v0),
    .vert0_valid_o         (valid_52_to_62_v0),
    .vert0_ready_i         (ready_62_to_52_v0),
    .vert1_data_i          (data_42_to_52_v1),
    .vert1_valid_i         (valid_42_to_52_v1),
    .vert1_ready_o         (ready_52_to_42_v1),
    .vert1_data_o          (data_52_to_62_v1),
    .vert1_valid_o         (valid_52_to_62_v1),
    .vert1_ready_i         (ready_62_to_52_v1),
    .local_data_i          (data_i[2][5]),
    .local_valid_i         (valid_i[2][5]),
    .local_ready_o         (ready_o[2][5]),
    .local_data_o          (data_o[2][5]),
    .local_valid_o         (valid_o[2][5]),
    .local_ready_i         (ready_i[2][5]),
    .credit_upd            (credit_upd)
);

/*Router 2,6*/    
cast_router #(
    .isUBM_list            (isUBM_list_2_6),
    .isFC_list             (isFC_list_2_6),
    .FCdn_list             (FCdn_list_2_6),
    .FCpl_list             (FCpl_list_2_6),
    .rt_file_list          (cast_rt_file_list_2_6)
)router_2_6(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_61_to_62),
    .west_valid_i          (valid_61_to_62),
    .west_ready_o          (ready_62_to_61),
    .west_data_o           (data_62_to_61),
    .west_valid_o          (valid_62_to_61),
    .west_ready_i          (ready_61_to_62),
    .east_data_i           (data_63_to_62),
    .east_valid_i          (valid_63_to_62),
    .east_ready_o          (ready_62_to_63),
    .east_data_o           (data_62_to_63),
    .east_valid_o          (valid_62_to_63),
    .east_ready_i          (ready_63_to_62),
    .vert0_data_i          (data_52_to_62_v0),
    .vert0_valid_i         (valid_52_to_62_v0),
    .vert0_ready_o         (ready_62_to_52_v0),
    .vert0_data_o          (data_62_to_72_v0),
    .vert0_valid_o         (valid_62_to_72_v0),
    .vert0_ready_i         (ready_72_to_62_v0),
    .vert1_data_i          (data_52_to_62_v1),
    .vert1_valid_i         (valid_52_to_62_v1),
    .vert1_ready_o         (ready_62_to_52_v1),
    .vert1_data_o          (data_62_to_72_v1),
    .vert1_valid_o         (valid_62_to_72_v1),
    .vert1_ready_i         (ready_72_to_62_v1),
    .local_data_i          (data_i[2][6]),
    .local_valid_i         (valid_i[2][6]),
    .local_ready_o         (ready_o[2][6]),
    .local_data_o          (data_o[2][6]),
    .local_valid_o         (valid_o[2][6]),
    .local_ready_i         (ready_i[2][6]),
    .credit_upd            (credit_upd)
);

/*Router 2,7*/    
cast_router #(
    .isUBM_list            (isUBM_list_2_7),
    .isFC_list             (isFC_list_2_7),
    .FCdn_list             (FCdn_list_2_7),
    .FCpl_list             (FCpl_list_2_7),
    .rt_file_list          (cast_rt_file_list_2_7)
)router_2_7(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_71_to_72),
    .west_valid_i          (valid_71_to_72),
    .west_ready_o          (ready_72_to_71),
    .west_data_o           (data_72_to_71),
    .west_valid_o          (valid_72_to_71),
    .west_ready_i          (ready_71_to_72),
    .east_data_i           (data_73_to_72),
    .east_valid_i          (valid_73_to_72),
    .east_ready_o          (ready_72_to_73),
    .east_data_o           (data_72_to_73),
    .east_valid_o          (valid_72_to_73),
    .east_ready_i          (ready_73_to_72),
    .vert0_data_i          (data_62_to_72_v0),
    .vert0_valid_i         (valid_62_to_72_v0),
    .vert0_ready_o         (ready_72_to_62_v0),
    .vert0_data_o          (data_72_to_82_v0),
    .vert0_valid_o         (valid_72_to_82_v0),
    .vert0_ready_i         (ready_82_to_72_v0),
    .vert1_data_i          (data_62_to_72_v1),
    .vert1_valid_i         (valid_62_to_72_v1),
    .vert1_ready_o         (ready_72_to_62_v1),
    .vert1_data_o          (data_72_to_82_v1),
    .vert1_valid_o         (valid_72_to_82_v1),
    .vert1_ready_i         (ready_82_to_72_v1),
    .local_data_i          (data_i[2][7]),
    .local_valid_i         (valid_i[2][7]),
    .local_ready_o         (ready_o[2][7]),
    .local_data_o          (data_o[2][7]),
    .local_valid_o         (valid_o[2][7]),
    .local_ready_i         (ready_i[2][7]),
    .credit_upd            (credit_upd)
);

/*Router 2,8*/    
cast_router #(
    .isUBM_list            (isUBM_list_2_8),
    .isFC_list             (isFC_list_2_8),
    .FCdn_list             (FCdn_list_2_8),
    .FCpl_list             (FCpl_list_2_8),
    .rt_file_list          (cast_rt_file_list_2_8)
)router_2_8(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_81_to_82),
    .west_valid_i          (valid_81_to_82),
    .west_ready_o          (ready_82_to_81),
    .west_data_o           (data_82_to_81),
    .west_valid_o          (valid_82_to_81),
    .west_ready_i          (ready_81_to_82),
    .east_data_i           (data_83_to_82),
    .east_valid_i          (valid_83_to_82),
    .east_ready_o          (ready_82_to_83),
    .east_data_o           (data_82_to_83),
    .east_valid_o          (valid_82_to_83),
    .east_ready_i          (ready_83_to_82),
    .vert0_data_i          (data_72_to_82_v0),
    .vert0_valid_i         (valid_72_to_82_v0),
    .vert0_ready_o         (ready_82_to_72_v0),
    .vert0_data_o          (data_82_to_92_v0),
    .vert0_valid_o         (valid_82_to_92_v0),
    .vert0_ready_i         (ready_92_to_82_v0),
    .vert1_data_i          (data_72_to_82_v1),
    .vert1_valid_i         (valid_72_to_82_v1),
    .vert1_ready_o         (ready_82_to_72_v1),
    .vert1_data_o          (data_82_to_92_v1),
    .vert1_valid_o         (valid_82_to_92_v1),
    .vert1_ready_i         (ready_92_to_82_v1),
    .local_data_i          (data_i[2][8]),
    .local_valid_i         (valid_i[2][8]),
    .local_ready_o         (ready_o[2][8]),
    .local_data_o          (data_o[2][8]),
    .local_valid_o         (valid_o[2][8]),
    .local_ready_i         (ready_i[2][8]),
    .credit_upd            (credit_upd)
);

/*Router 2,9*/    
cast_router #(
    .isUBM_list            (isUBM_list_2_9),
    .isFC_list             (isFC_list_2_9),
    .FCdn_list             (FCdn_list_2_9),
    .FCpl_list             (FCpl_list_2_9),
    .rt_file_list          (cast_rt_file_list_2_9)
)router_2_9(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_91_to_92),
    .west_valid_i          (valid_91_to_92),
    .west_ready_o          (ready_92_to_91),
    .west_data_o           (data_92_to_91),
    .west_valid_o          (valid_92_to_91),
    .west_ready_i          (ready_91_to_92),
    .east_data_i           (data_93_to_92),
    .east_valid_i          (valid_93_to_92),
    .east_ready_o          (ready_92_to_93),
    .east_data_o           (data_92_to_93),
    .east_valid_o          (valid_92_to_93),
    .east_ready_i          (ready_93_to_92),
    .vert0_data_i          (data_82_to_92_v0),
    .vert0_valid_i         (valid_82_to_92_v0),
    .vert0_ready_o         (ready_92_to_82_v0),
    .vert0_data_o          (data_92_to_102_v0),
    .vert0_valid_o         (valid_92_to_102_v0),
    .vert0_ready_i         (ready_102_to_92_v0),
    .vert1_data_i          (data_82_to_92_v1),
    .vert1_valid_i         (valid_82_to_92_v1),
    .vert1_ready_o         (ready_92_to_82_v1),
    .vert1_data_o          (data_92_to_102_v1),
    .vert1_valid_o         (valid_92_to_102_v1),
    .vert1_ready_i         (ready_102_to_92_v1),
    .local_data_i          (data_i[2][9]),
    .local_valid_i         (valid_i[2][9]),
    .local_ready_o         (ready_o[2][9]),
    .local_data_o          (data_o[2][9]),
    .local_valid_o         (valid_o[2][9]),
    .local_ready_i         (ready_i[2][9]),
    .credit_upd            (credit_upd)
);

/*Router 2,10*/    
cast_router #(
    .isUBM_list            (isUBM_list_2_10),
    .isFC_list             (isFC_list_2_10),
    .FCdn_list             (FCdn_list_2_10),
    .FCpl_list             (FCpl_list_2_10),
    .rt_file_list          (cast_rt_file_list_2_10)
)router_2_10(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_101_to_102),
    .west_valid_i          (valid_101_to_102),
    .west_ready_o          (ready_102_to_101),
    .west_data_o           (data_102_to_101),
    .west_valid_o          (valid_102_to_101),
    .west_ready_i          (ready_101_to_102),
    .east_data_i           (data_103_to_102),
    .east_valid_i          (valid_103_to_102),
    .east_ready_o          (ready_102_to_103),
    .east_data_o           (data_102_to_103),
    .east_valid_o          (valid_102_to_103),
    .east_ready_i          (ready_103_to_102),
    .vert0_data_i          (data_92_to_102_v0),
    .vert0_valid_i         (valid_92_to_102_v0),
    .vert0_ready_o         (ready_102_to_92_v0),
    .vert0_data_o          (data_102_to_112_v0),
    .vert0_valid_o         (valid_102_to_112_v0),
    .vert0_ready_i         (ready_112_to_102_v0),
    .vert1_data_i          (data_92_to_102_v1),
    .vert1_valid_i         (valid_92_to_102_v1),
    .vert1_ready_o         (ready_102_to_92_v1),
    .vert1_data_o          (data_102_to_112_v1),
    .vert1_valid_o         (valid_102_to_112_v1),
    .vert1_ready_i         (ready_112_to_102_v1),
    .local_data_i          (data_i[2][10]),
    .local_valid_i         (valid_i[2][10]),
    .local_ready_o         (ready_o[2][10]),
    .local_data_o          (data_o[2][10]),
    .local_valid_o         (valid_o[2][10]),
    .local_ready_i         (ready_i[2][10]),
    .credit_upd            (credit_upd)
);

/*Router 2,11*/    
cast_router #(
    .isUBM_list            (isUBM_list_2_11),
    .isFC_list             (isFC_list_2_11),
    .FCdn_list             (FCdn_list_2_11),
    .FCpl_list             (FCpl_list_2_11),
    .rt_file_list          (cast_rt_file_list_2_11)
)router_2_11(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_111_to_112),
    .west_valid_i          (valid_111_to_112),
    .west_ready_o          (ready_112_to_111),
    .west_data_o           (data_112_to_111),
    .west_valid_o          (valid_112_to_111),
    .west_ready_i          (ready_111_to_112),
    .east_data_i           (data_113_to_112),
    .east_valid_i          (valid_113_to_112),
    .east_ready_o          (ready_112_to_113),
    .east_data_o           (data_112_to_113),
    .east_valid_o          (valid_112_to_113),
    .east_ready_i          (ready_113_to_112),
    .vert0_data_i          (data_102_to_112_v0),
    .vert0_valid_i         (valid_102_to_112_v0),
    .vert0_ready_o         (ready_112_to_102_v0),
    .vert0_data_o          (data_112_to_122_v0),
    .vert0_valid_o         (valid_112_to_122_v0),
    .vert0_ready_i         (ready_122_to_112_v0),
    .vert1_data_i          (data_102_to_112_v1),
    .vert1_valid_i         (valid_102_to_112_v1),
    .vert1_ready_o         (ready_112_to_102_v1),
    .vert1_data_o          (data_112_to_122_v1),
    .vert1_valid_o         (valid_112_to_122_v1),
    .vert1_ready_i         (ready_122_to_112_v1),
    .local_data_i          (data_i[2][11]),
    .local_valid_i         (valid_i[2][11]),
    .local_ready_o         (ready_o[2][11]),
    .local_data_o          (data_o[2][11]),
    .local_valid_o         (valid_o[2][11]),
    .local_ready_i         (ready_i[2][11]),
    .credit_upd            (credit_upd)
);

/*Router 2,12*/    
cast_router #(
    .isUBM_list            (isUBM_list_2_12),
    .isFC_list             (isFC_list_2_12),
    .FCdn_list             (FCdn_list_2_12),
    .FCpl_list             (FCpl_list_2_12),
    .rt_file_list          (cast_rt_file_list_2_12)
)router_2_12(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_121_to_122),
    .west_valid_i          (valid_121_to_122),
    .west_ready_o          (ready_122_to_121),
    .west_data_o           (data_122_to_121),
    .west_valid_o          (valid_122_to_121),
    .west_ready_i          (ready_121_to_122),
    .east_data_i           (data_123_to_122),
    .east_valid_i          (valid_123_to_122),
    .east_ready_o          (ready_122_to_123),
    .east_data_o           (data_122_to_123),
    .east_valid_o          (valid_122_to_123),
    .east_ready_i          (ready_123_to_122),
    .vert0_data_i          (data_112_to_122_v0),
    .vert0_valid_i         (valid_112_to_122_v0),
    .vert0_ready_o         (ready_122_to_112_v0),
    .vert0_data_o          (data_122_to_132_v0),
    .vert0_valid_o         (valid_122_to_132_v0),
    .vert0_ready_i         (ready_132_to_122_v0),
    .vert1_data_i          (data_112_to_122_v1),
    .vert1_valid_i         (valid_112_to_122_v1),
    .vert1_ready_o         (ready_122_to_112_v1),
    .vert1_data_o          (data_122_to_132_v1),
    .vert1_valid_o         (valid_122_to_132_v1),
    .vert1_ready_i         (ready_132_to_122_v1),
    .local_data_i          (data_i[2][12]),
    .local_valid_i         (valid_i[2][12]),
    .local_ready_o         (ready_o[2][12]),
    .local_data_o          (data_o[2][12]),
    .local_valid_o         (valid_o[2][12]),
    .local_ready_i         (ready_i[2][12]),
    .credit_upd            (credit_upd)
);

/*Router 2,13*/    
cast_router #(
    .isUBM_list            (isUBM_list_2_13),
    .isFC_list             (isFC_list_2_13),
    .FCdn_list             (FCdn_list_2_13),
    .FCpl_list             (FCpl_list_2_13),
    .rt_file_list          (cast_rt_file_list_2_13)
)router_2_13(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_131_to_132),
    .west_valid_i          (valid_131_to_132),
    .west_ready_o          (ready_132_to_131),
    .west_data_o           (data_132_to_131),
    .west_valid_o          (valid_132_to_131),
    .west_ready_i          (ready_131_to_132),
    .east_data_i           (data_133_to_132),
    .east_valid_i          (valid_133_to_132),
    .east_ready_o          (ready_132_to_133),
    .east_data_o           (data_132_to_133),
    .east_valid_o          (valid_132_to_133),
    .east_ready_i          (ready_133_to_132),
    .vert0_data_i          (data_122_to_132_v0),
    .vert0_valid_i         (valid_122_to_132_v0),
    .vert0_ready_o         (ready_132_to_122_v0),
    .vert0_data_o          (data_132_to_142_v0),
    .vert0_valid_o         (valid_132_to_142_v0),
    .vert0_ready_i         (ready_142_to_132_v0),
    .vert1_data_i          (data_122_to_132_v1),
    .vert1_valid_i         (valid_122_to_132_v1),
    .vert1_ready_o         (ready_132_to_122_v1),
    .vert1_data_o          (data_132_to_142_v1),
    .vert1_valid_o         (valid_132_to_142_v1),
    .vert1_ready_i         (ready_142_to_132_v1),
    .local_data_i          (data_i[2][13]),
    .local_valid_i         (valid_i[2][13]),
    .local_ready_o         (ready_o[2][13]),
    .local_data_o          (data_o[2][13]),
    .local_valid_o         (valid_o[2][13]),
    .local_ready_i         (ready_i[2][13]),
    .credit_upd            (credit_upd)
);

/*Router 2,14*/    
cast_router #(
    .isUBM_list            (isUBM_list_2_14),
    .isFC_list             (isFC_list_2_14),
    .FCdn_list             (FCdn_list_2_14),
    .FCpl_list             (FCpl_list_2_14),
    .rt_file_list          (cast_rt_file_list_2_14)
)router_2_14(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_141_to_142),
    .west_valid_i          (valid_141_to_142),
    .west_ready_o          (ready_142_to_141),
    .west_data_o           (data_142_to_141),
    .west_valid_o          (valid_142_to_141),
    .west_ready_i          (ready_141_to_142),
    .east_data_i           (data_143_to_142),
    .east_valid_i          (valid_143_to_142),
    .east_ready_o          (ready_142_to_143),
    .east_data_o           (data_142_to_143),
    .east_valid_o          (valid_142_to_143),
    .east_ready_i          (ready_143_to_142),
    .vert0_data_i          (data_132_to_142_v0),
    .vert0_valid_i         (valid_132_to_142_v0),
    .vert0_ready_o         (ready_142_to_132_v0),
    .vert0_data_o          (data_142_to_152_v0),
    .vert0_valid_o         (valid_142_to_152_v0),
    .vert0_ready_i         (ready_152_to_142_v0),
    .vert1_data_i          (data_132_to_142_v1),
    .vert1_valid_i         (valid_132_to_142_v1),
    .vert1_ready_o         (ready_142_to_132_v1),
    .vert1_data_o          (data_142_to_152_v1),
    .vert1_valid_o         (valid_142_to_152_v1),
    .vert1_ready_i         (ready_152_to_142_v1),
    .local_data_i          (data_i[2][14]),
    .local_valid_i         (valid_i[2][14]),
    .local_ready_o         (ready_o[2][14]),
    .local_data_o          (data_o[2][14]),
    .local_valid_o         (valid_o[2][14]),
    .local_ready_i         (ready_i[2][14]),
    .credit_upd            (credit_upd)
);

/*Router 2,15*/    
cast_router #(
    .isUBM_list            (isUBM_list_2_15),
    .isFC_list             (isFC_list_2_15),
    .FCdn_list             (FCdn_list_2_15),
    .FCpl_list             (FCpl_list_2_15),
    .rt_file_list          (cast_rt_file_list_2_15)
)router_2_15(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_151_to_152),
    .west_valid_i          (valid_151_to_152),
    .west_ready_o          (ready_152_to_151),
    .west_data_o           (data_152_to_151),
    .west_valid_o          (valid_152_to_151),
    .west_ready_i          (ready_151_to_152),
    .east_data_i           (data_153_to_152),
    .east_valid_i          (valid_153_to_152),
    .east_ready_o          (ready_152_to_153),
    .east_data_o           (data_152_to_153),
    .east_valid_o          (valid_152_to_153),
    .east_ready_i          (ready_153_to_152),
    .vert0_data_i          (data_142_to_152_v0),
    .vert0_valid_i         (valid_142_to_152_v0),
    .vert0_ready_o         (ready_152_to_142_v0),
    .vert0_data_o          (data_152_to_162_v0),
    .vert0_valid_o         (valid_152_to_162_v0),
    .vert0_ready_i         (ready_162_to_152_v0),
    .vert1_data_i          (data_142_to_152_v1),
    .vert1_valid_i         (valid_142_to_152_v1),
    .vert1_ready_o         (ready_152_to_142_v1),
    .vert1_data_o          (data_152_to_162_v1),
    .vert1_valid_o         (valid_152_to_162_v1),
    .vert1_ready_i         (ready_162_to_152_v1),
    .local_data_i          (data_i[2][15]),
    .local_valid_i         (valid_i[2][15]),
    .local_ready_o         (ready_o[2][15]),
    .local_data_o          (data_o[2][15]),
    .local_valid_o         (valid_o[2][15]),
    .local_ready_i         (ready_i[2][15]),
    .credit_upd            (credit_upd)
);

/*Router 2,16*/    
cast_router #(
    .isUBM_list            (isUBM_list_2_16),
    .isFC_list             (isFC_list_2_16),
    .FCdn_list             (FCdn_list_2_16),
    .FCpl_list             (FCpl_list_2_16),
    .rt_file_list          (cast_rt_file_list_2_16)
)router_2_16(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_161_to_162),
    .west_valid_i          (valid_161_to_162),
    .west_ready_o          (ready_162_to_161),
    .west_data_o           (data_162_to_161),
    .west_valid_o          (valid_162_to_161),
    .west_ready_i          (ready_161_to_162),
    .east_data_i           (data_163_to_162),
    .east_valid_i          (valid_163_to_162),
    .east_ready_o          (ready_162_to_163),
    .east_data_o           (data_162_to_163),
    .east_valid_o          (valid_162_to_163),
    .east_ready_i          (ready_163_to_162),
    .vert0_data_i          (data_152_to_162_v0),
    .vert0_valid_i         (valid_152_to_162_v0),
    .vert0_ready_o         (ready_162_to_152_v0),
    .vert0_data_o          (data_162_to_172_v0),
    .vert0_valid_o         (valid_162_to_172_v0),
    .vert0_ready_i         (ready_172_to_162_v0),
    .vert1_data_i          (data_152_to_162_v1),
    .vert1_valid_i         (valid_152_to_162_v1),
    .vert1_ready_o         (ready_162_to_152_v1),
    .vert1_data_o          (data_162_to_172_v1),
    .vert1_valid_o         (valid_162_to_172_v1),
    .vert1_ready_i         (ready_172_to_162_v1),
    .local_data_i          (data_i[2][16]),
    .local_valid_i         (valid_i[2][16]),
    .local_ready_o         (ready_o[2][16]),
    .local_data_o          (data_o[2][16]),
    .local_valid_o         (valid_o[2][16]),
    .local_ready_i         (ready_i[2][16]),
    .credit_upd            (credit_upd)
);

/*Router 2,17*/    
cast_router #(
    .isUBM_list            (isUBM_list_2_17),
    .isFC_list             (isFC_list_2_17),
    .FCdn_list             (FCdn_list_2_17),
    .FCpl_list             (FCpl_list_2_17),
    .rt_file_list          (cast_rt_file_list_2_17)
)router_2_17(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_171_to_172),
    .west_valid_i          (valid_171_to_172),
    .west_ready_o          (ready_172_to_171),
    .west_data_o           (data_172_to_171),
    .west_valid_o          (valid_172_to_171),
    .west_ready_i          (ready_171_to_172),
    .east_data_i           (data_173_to_172),
    .east_valid_i          (valid_173_to_172),
    .east_ready_o          (ready_172_to_173),
    .east_data_o           (data_172_to_173),
    .east_valid_o          (valid_172_to_173),
    .east_ready_i          (ready_173_to_172),
    .vert0_data_i          (data_162_to_172_v0),
    .vert0_valid_i         (valid_162_to_172_v0),
    .vert0_ready_o         (ready_172_to_162_v0),
    .vert0_data_o          (data_172_to_182_v0),
    .vert0_valid_o         (valid_172_to_182_v0),
    .vert0_ready_i         (ready_182_to_172_v0),
    .vert1_data_i          (data_162_to_172_v1),
    .vert1_valid_i         (valid_162_to_172_v1),
    .vert1_ready_o         (ready_172_to_162_v1),
    .vert1_data_o          (data_172_to_182_v1),
    .vert1_valid_o         (valid_172_to_182_v1),
    .vert1_ready_i         (ready_182_to_172_v1),
    .local_data_i          (data_i[2][17]),
    .local_valid_i         (valid_i[2][17]),
    .local_ready_o         (ready_o[2][17]),
    .local_data_o          (data_o[2][17]),
    .local_valid_o         (valid_o[2][17]),
    .local_ready_i         (ready_i[2][17]),
    .credit_upd            (credit_upd)
);

/*Router 2,18*/    
cast_router #(
    .isUBM_list            (isUBM_list_2_18),
    .isFC_list             (isFC_list_2_18),
    .FCdn_list             (FCdn_list_2_18),
    .FCpl_list             (FCpl_list_2_18),
    .rt_file_list          (cast_rt_file_list_2_18)
)router_2_18(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_181_to_182),
    .west_valid_i          (valid_181_to_182),
    .west_ready_o          (ready_182_to_181),
    .west_data_o           (data_182_to_181),
    .west_valid_o          (valid_182_to_181),
    .west_ready_i          (ready_181_to_182),
    .east_data_i           (data_183_to_182),
    .east_valid_i          (valid_183_to_182),
    .east_ready_o          (ready_182_to_183),
    .east_data_o           (data_182_to_183),
    .east_valid_o          (valid_182_to_183),
    .east_ready_i          (ready_183_to_182),
    .vert0_data_i          (data_172_to_182_v0),
    .vert0_valid_i         (valid_172_to_182_v0),
    .vert0_ready_o         (ready_182_to_172_v0),
    .vert0_data_o          (data_182_to_192_v0),
    .vert0_valid_o         (valid_182_to_192_v0),
    .vert0_ready_i         (ready_192_to_182_v0),
    .vert1_data_i          (data_172_to_182_v1),
    .vert1_valid_i         (valid_172_to_182_v1),
    .vert1_ready_o         (ready_182_to_172_v1),
    .vert1_data_o          (data_182_to_192_v1),
    .vert1_valid_o         (valid_182_to_192_v1),
    .vert1_ready_i         (ready_192_to_182_v1),
    .local_data_i          (data_i[2][18]),
    .local_valid_i         (valid_i[2][18]),
    .local_ready_o         (ready_o[2][18]),
    .local_data_o          (data_o[2][18]),
    .local_valid_o         (valid_o[2][18]),
    .local_ready_i         (ready_i[2][18]),
    .credit_upd            (credit_upd)
);

/*Router 2,19*/    
cast_router #(
    .isUBM_list            (isUBM_list_2_19),
    .isFC_list             (isFC_list_2_19),
    .FCdn_list             (FCdn_list_2_19),
    .FCpl_list             (FCpl_list_2_19),
    .rt_file_list          (cast_rt_file_list_2_19)
)router_2_19(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_191_to_192),
    .west_valid_i          (valid_191_to_192),
    .west_ready_o          (ready_192_to_191),
    .west_data_o           (data_192_to_191),
    .west_valid_o          (valid_192_to_191),
    .west_ready_i          (ready_191_to_192),
    .east_data_i           (data_193_to_192),
    .east_valid_i          (valid_193_to_192),
    .east_ready_o          (ready_192_to_193),
    .east_data_o           (data_192_to_193),
    .east_valid_o          (valid_192_to_193),
    .east_ready_i          (ready_193_to_192),
    .vert0_data_i          (data_182_to_192_v0),
    .vert0_valid_i         (valid_182_to_192_v0),
    .vert0_ready_o         (ready_192_to_182_v0),
    .vert0_data_o          (data_192_to_202_v0),
    .vert0_valid_o         (valid_192_to_202_v0),
    .vert0_ready_i         (ready_202_to_192_v0),
    .vert1_data_i          (data_182_to_192_v1),
    .vert1_valid_i         (valid_182_to_192_v1),
    .vert1_ready_o         (ready_192_to_182_v1),
    .vert1_data_o          (data_192_to_202_v1),
    .vert1_valid_o         (valid_192_to_202_v1),
    .vert1_ready_i         (ready_202_to_192_v1),
    .local_data_i          (data_i[2][19]),
    .local_valid_i         (valid_i[2][19]),
    .local_ready_o         (ready_o[2][19]),
    .local_data_o          (data_o[2][19]),
    .local_valid_o         (valid_o[2][19]),
    .local_ready_i         (ready_i[2][19]),
    .credit_upd            (credit_upd)
);

/*Router 2,20*/    
cast_router #(
    .isUBM_list            (isUBM_list_2_20),
    .isFC_list             (isFC_list_2_20),
    .FCdn_list             (FCdn_list_2_20),
    .FCpl_list             (FCpl_list_2_20),
    .rt_file_list          (cast_rt_file_list_2_20)
)router_2_20(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_201_to_202),
    .west_valid_i          (valid_201_to_202),
    .west_ready_o          (ready_202_to_201),
    .west_data_o           (data_202_to_201),
    .west_valid_o          (valid_202_to_201),
    .west_ready_i          (ready_201_to_202),
    .east_data_i           (data_203_to_202),
    .east_valid_i          (valid_203_to_202),
    .east_ready_o          (ready_202_to_203),
    .east_data_o           (data_202_to_203),
    .east_valid_o          (valid_202_to_203),
    .east_ready_i          (ready_203_to_202),
    .vert0_data_i          (data_192_to_202_v0),
    .vert0_valid_i         (valid_192_to_202_v0),
    .vert0_ready_o         (ready_202_to_192_v0),
    .vert0_data_o          (data_202_to_212_v0),
    .vert0_valid_o         (valid_202_to_212_v0),
    .vert0_ready_i         (ready_212_to_202_v0),
    .vert1_data_i          (data_192_to_202_v1),
    .vert1_valid_i         (valid_192_to_202_v1),
    .vert1_ready_o         (ready_202_to_192_v1),
    .vert1_data_o          (data_202_to_212_v1),
    .vert1_valid_o         (valid_202_to_212_v1),
    .vert1_ready_i         (ready_212_to_202_v1),
    .local_data_i          (data_i[2][20]),
    .local_valid_i         (valid_i[2][20]),
    .local_ready_o         (ready_o[2][20]),
    .local_data_o          (data_o[2][20]),
    .local_valid_o         (valid_o[2][20]),
    .local_ready_i         (ready_i[2][20]),
    .credit_upd            (credit_upd)
);

/*Router 2,21*/    
cast_router #(
    .isUBM_list            (isUBM_list_2_21),
    .isFC_list             (isFC_list_2_21),
    .FCdn_list             (FCdn_list_2_21),
    .FCpl_list             (FCpl_list_2_21),
    .rt_file_list          (cast_rt_file_list_2_21)
)router_2_21(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_211_to_212),
    .west_valid_i          (valid_211_to_212),
    .west_ready_o          (ready_212_to_211),
    .west_data_o           (data_212_to_211),
    .west_valid_o          (valid_212_to_211),
    .west_ready_i          (ready_211_to_212),
    .east_data_i           (data_213_to_212),
    .east_valid_i          (valid_213_to_212),
    .east_ready_o          (ready_212_to_213),
    .east_data_o           (data_212_to_213),
    .east_valid_o          (valid_212_to_213),
    .east_ready_i          (ready_213_to_212),
    .vert0_data_i          (data_202_to_212_v0),
    .vert0_valid_i         (valid_202_to_212_v0),
    .vert0_ready_o         (ready_212_to_202_v0),
    .vert0_data_o          (data_212_to_222_v0),
    .vert0_valid_o         (valid_212_to_222_v0),
    .vert0_ready_i         (ready_222_to_212_v0),
    .vert1_data_i          (data_202_to_212_v1),
    .vert1_valid_i         (valid_202_to_212_v1),
    .vert1_ready_o         (ready_212_to_202_v1),
    .vert1_data_o          (data_212_to_222_v1),
    .vert1_valid_o         (valid_212_to_222_v1),
    .vert1_ready_i         (ready_222_to_212_v1),
    .local_data_i          (data_i[2][21]),
    .local_valid_i         (valid_i[2][21]),
    .local_ready_o         (ready_o[2][21]),
    .local_data_o          (data_o[2][21]),
    .local_valid_o         (valid_o[2][21]),
    .local_ready_i         (ready_i[2][21]),
    .credit_upd            (credit_upd)
);

/*Router 2,22*/    
cast_router #(
    .isUBM_list            (isUBM_list_2_22),
    .isFC_list             (isFC_list_2_22),
    .FCdn_list             (FCdn_list_2_22),
    .FCpl_list             (FCpl_list_2_22),
    .rt_file_list          (cast_rt_file_list_2_22)
)router_2_22(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_221_to_222),
    .west_valid_i          (valid_221_to_222),
    .west_ready_o          (ready_222_to_221),
    .west_data_o           (data_222_to_221),
    .west_valid_o          (valid_222_to_221),
    .west_ready_i          (ready_221_to_222),
    .east_data_i           (data_223_to_222),
    .east_valid_i          (valid_223_to_222),
    .east_ready_o          (ready_222_to_223),
    .east_data_o           (data_222_to_223),
    .east_valid_o          (valid_222_to_223),
    .east_ready_i          (ready_223_to_222),
    .vert0_data_i          (data_212_to_222_v0),
    .vert0_valid_i         (valid_212_to_222_v0),
    .vert0_ready_o         (ready_222_to_212_v0),
    .vert0_data_o          (data_222_to_232_v0),
    .vert0_valid_o         (valid_222_to_232_v0),
    .vert0_ready_i         (ready_232_to_222_v0),
    .vert1_data_i          (data_212_to_222_v1),
    .vert1_valid_i         (valid_212_to_222_v1),
    .vert1_ready_o         (ready_222_to_212_v1),
    .vert1_data_o          (data_222_to_232_v1),
    .vert1_valid_o         (valid_222_to_232_v1),
    .vert1_ready_i         (ready_232_to_222_v1),
    .local_data_i          (data_i[2][22]),
    .local_valid_i         (valid_i[2][22]),
    .local_ready_o         (ready_o[2][22]),
    .local_data_o          (data_o[2][22]),
    .local_valid_o         (valid_o[2][22]),
    .local_ready_i         (ready_i[2][22]),
    .credit_upd            (credit_upd)
);

/*Router 2,23*/    
cast_router #(
    .isUBM_list            (isUBM_list_2_23),
    .isFC_list             (isFC_list_2_23),
    .FCdn_list             (FCdn_list_2_23),
    .FCpl_list             (FCpl_list_2_23),
    .rt_file_list          (cast_rt_file_list_2_23)
)router_2_23(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_231_to_232),
    .west_valid_i          (valid_231_to_232),
    .west_ready_o          (ready_232_to_231),
    .west_data_o           (data_232_to_231),
    .west_valid_o          (valid_232_to_231),
    .west_ready_i          (ready_231_to_232),
    .east_data_i           (data_233_to_232),
    .east_valid_i          (valid_233_to_232),
    .east_ready_o          (ready_232_to_233),
    .east_data_o           (data_232_to_233),
    .east_valid_o          (valid_232_to_233),
    .east_ready_i          (ready_233_to_232),
    .vert0_data_i          (data_222_to_232_v0),
    .vert0_valid_i         (valid_222_to_232_v0),
    .vert0_ready_o         (ready_232_to_222_v0),
    .vert0_data_o          (data_232_to_242_v0),
    .vert0_valid_o         (valid_232_to_242_v0),
    .vert0_ready_i         (ready_242_to_232_v0),
    .vert1_data_i          (data_222_to_232_v1),
    .vert1_valid_i         (valid_222_to_232_v1),
    .vert1_ready_o         (ready_232_to_222_v1),
    .vert1_data_o          (data_232_to_242_v1),
    .vert1_valid_o         (valid_232_to_242_v1),
    .vert1_ready_i         (ready_242_to_232_v1),
    .local_data_i          (data_i[2][23]),
    .local_valid_i         (valid_i[2][23]),
    .local_ready_o         (ready_o[2][23]),
    .local_data_o          (data_o[2][23]),
    .local_valid_o         (valid_o[2][23]),
    .local_ready_i         (ready_i[2][23]),
    .credit_upd            (credit_upd)
);

/*Router 2,24*/    
cast_router #(
    .isUBM_list            (isUBM_list_2_24),
    .isFC_list             (isFC_list_2_24),
    .FCdn_list             (FCdn_list_2_24),
    .FCpl_list             (FCpl_list_2_24),
    .rt_file_list          (cast_rt_file_list_2_24)
)router_2_24(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_241_to_242),
    .west_valid_i          (valid_241_to_242),
    .west_ready_o          (ready_242_to_241),
    .west_data_o           (data_242_to_241),
    .west_valid_o          (valid_242_to_241),
    .west_ready_i          (ready_241_to_242),
    .east_data_i           (data_243_to_242),
    .east_valid_i          (valid_243_to_242),
    .east_ready_o          (ready_242_to_243),
    .east_data_o           (data_242_to_243),
    .east_valid_o          (valid_242_to_243),
    .east_ready_i          (ready_243_to_242),
    .vert0_data_i          (data_232_to_242_v0),
    .vert0_valid_i         (valid_232_to_242_v0),
    .vert0_ready_o         (ready_242_to_232_v0),
    .vert0_data_o          (),
    .vert0_valid_o         (),
    .vert0_ready_i         (1'b0),
    .vert1_data_i          (data_232_to_242_v1),
    .vert1_valid_i         (valid_232_to_242_v1),
    .vert1_ready_o         (ready_242_to_232_v1),
    .vert1_data_o          (),
    .vert1_valid_o         (),
    .vert1_ready_i         (1'b0),
    .local_data_i          (data_i[2][24]),
    .local_valid_i         (valid_i[2][24]),
    .local_ready_o         (ready_o[2][24]),
    .local_data_o          (data_o[2][24]),
    .local_valid_o         (valid_o[2][24]),
    .local_ready_i         (ready_i[2][24]),
    .credit_upd            (credit_upd)
);

/*Router 3,0*/    
cast_router #(
    .isUBM_list            (isUBM_list_3_0),
    .isFC_list             (isFC_list_3_0),
    .FCdn_list             (FCdn_list_3_0),
    .FCpl_list             (FCpl_list_3_0),
    .rt_file_list          (cast_rt_file_list_3_0)
)router_3_0(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_2_to_3),
    .west_valid_i          (valid_2_to_3),
    .west_ready_o          (ready_3_to_2),
    .west_data_o           (data_3_to_2),
    .west_valid_o          (valid_3_to_2),
    .west_ready_i          (ready_2_to_3),
    .east_data_i           (data_4_to_3),
    .east_valid_i          (valid_4_to_3),
    .east_ready_o          (ready_3_to_4),
    .east_data_o           (data_3_to_4),
    .east_valid_o          (valid_3_to_4),
    .east_ready_i          (ready_4_to_3),
    .vert0_data_i          (34'b0),
    .vert0_valid_i         (1'b0),
    .vert0_ready_o         (),
    .vert0_data_o          (data_3_to_13_v0),
    .vert0_valid_o         (valid_3_to_13_v0),
    .vert0_ready_i         (ready_13_to_3_v0),
    .vert1_data_i          (34'b0),
    .vert1_valid_i         (1'b0),
    .vert1_ready_o         (),
    .vert1_data_o          (data_3_to_13_v1),
    .vert1_valid_o         (valid_3_to_13_v1),
    .vert1_ready_i         (ready_13_to_3_v1),
    .local_data_i          (data_i[3][0]),
    .local_valid_i         (valid_i[3][0]),
    .local_ready_o         (ready_o[3][0]),
    .local_data_o          (data_o[3][0]),
    .local_valid_o         (valid_o[3][0]),
    .local_ready_i         (ready_i[3][0]),
    .credit_upd            (credit_upd)
);

/*Router 3,1*/    
cast_router #(
    .isUBM_list            (isUBM_list_3_1),
    .isFC_list             (isFC_list_3_1),
    .FCdn_list             (FCdn_list_3_1),
    .FCpl_list             (FCpl_list_3_1),
    .rt_file_list          (cast_rt_file_list_3_1)
)router_3_1(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_12_to_13),
    .west_valid_i          (valid_12_to_13),
    .west_ready_o          (ready_13_to_12),
    .west_data_o           (data_13_to_12),
    .west_valid_o          (valid_13_to_12),
    .west_ready_i          (ready_12_to_13),
    .east_data_i           (data_14_to_13),
    .east_valid_i          (valid_14_to_13),
    .east_ready_o          (ready_13_to_14),
    .east_data_o           (data_13_to_14),
    .east_valid_o          (valid_13_to_14),
    .east_ready_i          (ready_14_to_13),
    .vert0_data_i          (data_3_to_13_v0),
    .vert0_valid_i         (valid_3_to_13_v0),
    .vert0_ready_o         (ready_13_to_3_v0),
    .vert0_data_o          (data_13_to_23_v0),
    .vert0_valid_o         (valid_13_to_23_v0),
    .vert0_ready_i         (ready_23_to_13_v0),
    .vert1_data_i          (data_3_to_13_v1),
    .vert1_valid_i         (valid_3_to_13_v1),
    .vert1_ready_o         (ready_13_to_3_v1),
    .vert1_data_o          (data_13_to_23_v1),
    .vert1_valid_o         (valid_13_to_23_v1),
    .vert1_ready_i         (ready_23_to_13_v1),
    .local_data_i          (data_i[3][1]),
    .local_valid_i         (valid_i[3][1]),
    .local_ready_o         (ready_o[3][1]),
    .local_data_o          (data_o[3][1]),
    .local_valid_o         (valid_o[3][1]),
    .local_ready_i         (ready_i[3][1]),
    .credit_upd            (credit_upd)
);

/*Router 3,2*/    
cast_router #(
    .isUBM_list            (isUBM_list_3_2),
    .isFC_list             (isFC_list_3_2),
    .FCdn_list             (FCdn_list_3_2),
    .FCpl_list             (FCpl_list_3_2),
    .rt_file_list          (cast_rt_file_list_3_2)
)router_3_2(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_22_to_23),
    .west_valid_i          (valid_22_to_23),
    .west_ready_o          (ready_23_to_22),
    .west_data_o           (data_23_to_22),
    .west_valid_o          (valid_23_to_22),
    .west_ready_i          (ready_22_to_23),
    .east_data_i           (data_24_to_23),
    .east_valid_i          (valid_24_to_23),
    .east_ready_o          (ready_23_to_24),
    .east_data_o           (data_23_to_24),
    .east_valid_o          (valid_23_to_24),
    .east_ready_i          (ready_24_to_23),
    .vert0_data_i          (data_13_to_23_v0),
    .vert0_valid_i         (valid_13_to_23_v0),
    .vert0_ready_o         (ready_23_to_13_v0),
    .vert0_data_o          (data_23_to_33_v0),
    .vert0_valid_o         (valid_23_to_33_v0),
    .vert0_ready_i         (ready_33_to_23_v0),
    .vert1_data_i          (data_13_to_23_v1),
    .vert1_valid_i         (valid_13_to_23_v1),
    .vert1_ready_o         (ready_23_to_13_v1),
    .vert1_data_o          (data_23_to_33_v1),
    .vert1_valid_o         (valid_23_to_33_v1),
    .vert1_ready_i         (ready_33_to_23_v1),
    .local_data_i          (data_i[3][2]),
    .local_valid_i         (valid_i[3][2]),
    .local_ready_o         (ready_o[3][2]),
    .local_data_o          (data_o[3][2]),
    .local_valid_o         (valid_o[3][2]),
    .local_ready_i         (ready_i[3][2]),
    .credit_upd            (credit_upd)
);

/*Router 3,3*/    
cast_router #(
    .isUBM_list            (isUBM_list_3_3),
    .isFC_list             (isFC_list_3_3),
    .FCdn_list             (FCdn_list_3_3),
    .FCpl_list             (FCpl_list_3_3),
    .rt_file_list          (cast_rt_file_list_3_3)
)router_3_3(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_32_to_33),
    .west_valid_i          (valid_32_to_33),
    .west_ready_o          (ready_33_to_32),
    .west_data_o           (data_33_to_32),
    .west_valid_o          (valid_33_to_32),
    .west_ready_i          (ready_32_to_33),
    .east_data_i           (data_34_to_33),
    .east_valid_i          (valid_34_to_33),
    .east_ready_o          (ready_33_to_34),
    .east_data_o           (data_33_to_34),
    .east_valid_o          (valid_33_to_34),
    .east_ready_i          (ready_34_to_33),
    .vert0_data_i          (data_23_to_33_v0),
    .vert0_valid_i         (valid_23_to_33_v0),
    .vert0_ready_o         (ready_33_to_23_v0),
    .vert0_data_o          (data_33_to_43_v0),
    .vert0_valid_o         (valid_33_to_43_v0),
    .vert0_ready_i         (ready_43_to_33_v0),
    .vert1_data_i          (data_23_to_33_v1),
    .vert1_valid_i         (valid_23_to_33_v1),
    .vert1_ready_o         (ready_33_to_23_v1),
    .vert1_data_o          (data_33_to_43_v1),
    .vert1_valid_o         (valid_33_to_43_v1),
    .vert1_ready_i         (ready_43_to_33_v1),
    .local_data_i          (data_i[3][3]),
    .local_valid_i         (valid_i[3][3]),
    .local_ready_o         (ready_o[3][3]),
    .local_data_o          (data_o[3][3]),
    .local_valid_o         (valid_o[3][3]),
    .local_ready_i         (ready_i[3][3]),
    .credit_upd            (credit_upd)
);

/*Router 3,4*/    
cast_router #(
    .isUBM_list            (isUBM_list_3_4),
    .isFC_list             (isFC_list_3_4),
    .FCdn_list             (FCdn_list_3_4),
    .FCpl_list             (FCpl_list_3_4),
    .rt_file_list          (cast_rt_file_list_3_4)
)router_3_4(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_42_to_43),
    .west_valid_i          (valid_42_to_43),
    .west_ready_o          (ready_43_to_42),
    .west_data_o           (data_43_to_42),
    .west_valid_o          (valid_43_to_42),
    .west_ready_i          (ready_42_to_43),
    .east_data_i           (data_44_to_43),
    .east_valid_i          (valid_44_to_43),
    .east_ready_o          (ready_43_to_44),
    .east_data_o           (data_43_to_44),
    .east_valid_o          (valid_43_to_44),
    .east_ready_i          (ready_44_to_43),
    .vert0_data_i          (data_33_to_43_v0),
    .vert0_valid_i         (valid_33_to_43_v0),
    .vert0_ready_o         (ready_43_to_33_v0),
    .vert0_data_o          (data_43_to_53_v0),
    .vert0_valid_o         (valid_43_to_53_v0),
    .vert0_ready_i         (ready_53_to_43_v0),
    .vert1_data_i          (data_33_to_43_v1),
    .vert1_valid_i         (valid_33_to_43_v1),
    .vert1_ready_o         (ready_43_to_33_v1),
    .vert1_data_o          (data_43_to_53_v1),
    .vert1_valid_o         (valid_43_to_53_v1),
    .vert1_ready_i         (ready_53_to_43_v1),
    .local_data_i          (data_i[3][4]),
    .local_valid_i         (valid_i[3][4]),
    .local_ready_o         (ready_o[3][4]),
    .local_data_o          (data_o[3][4]),
    .local_valid_o         (valid_o[3][4]),
    .local_ready_i         (ready_i[3][4]),
    .credit_upd            (credit_upd)
);

/*Router 3,5*/    
cast_router #(
    .isUBM_list            (isUBM_list_3_5),
    .isFC_list             (isFC_list_3_5),
    .FCdn_list             (FCdn_list_3_5),
    .FCpl_list             (FCpl_list_3_5),
    .rt_file_list          (cast_rt_file_list_3_5)
)router_3_5(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_52_to_53),
    .west_valid_i          (valid_52_to_53),
    .west_ready_o          (ready_53_to_52),
    .west_data_o           (data_53_to_52),
    .west_valid_o          (valid_53_to_52),
    .west_ready_i          (ready_52_to_53),
    .east_data_i           (data_54_to_53),
    .east_valid_i          (valid_54_to_53),
    .east_ready_o          (ready_53_to_54),
    .east_data_o           (data_53_to_54),
    .east_valid_o          (valid_53_to_54),
    .east_ready_i          (ready_54_to_53),
    .vert0_data_i          (data_43_to_53_v0),
    .vert0_valid_i         (valid_43_to_53_v0),
    .vert0_ready_o         (ready_53_to_43_v0),
    .vert0_data_o          (data_53_to_63_v0),
    .vert0_valid_o         (valid_53_to_63_v0),
    .vert0_ready_i         (ready_63_to_53_v0),
    .vert1_data_i          (data_43_to_53_v1),
    .vert1_valid_i         (valid_43_to_53_v1),
    .vert1_ready_o         (ready_53_to_43_v1),
    .vert1_data_o          (data_53_to_63_v1),
    .vert1_valid_o         (valid_53_to_63_v1),
    .vert1_ready_i         (ready_63_to_53_v1),
    .local_data_i          (data_i[3][5]),
    .local_valid_i         (valid_i[3][5]),
    .local_ready_o         (ready_o[3][5]),
    .local_data_o          (data_o[3][5]),
    .local_valid_o         (valid_o[3][5]),
    .local_ready_i         (ready_i[3][5]),
    .credit_upd            (credit_upd)
);

/*Router 3,6*/    
cast_router #(
    .isUBM_list            (isUBM_list_3_6),
    .isFC_list             (isFC_list_3_6),
    .FCdn_list             (FCdn_list_3_6),
    .FCpl_list             (FCpl_list_3_6),
    .rt_file_list          (cast_rt_file_list_3_6)
)router_3_6(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_62_to_63),
    .west_valid_i          (valid_62_to_63),
    .west_ready_o          (ready_63_to_62),
    .west_data_o           (data_63_to_62),
    .west_valid_o          (valid_63_to_62),
    .west_ready_i          (ready_62_to_63),
    .east_data_i           (data_64_to_63),
    .east_valid_i          (valid_64_to_63),
    .east_ready_o          (ready_63_to_64),
    .east_data_o           (data_63_to_64),
    .east_valid_o          (valid_63_to_64),
    .east_ready_i          (ready_64_to_63),
    .vert0_data_i          (data_53_to_63_v0),
    .vert0_valid_i         (valid_53_to_63_v0),
    .vert0_ready_o         (ready_63_to_53_v0),
    .vert0_data_o          (data_63_to_73_v0),
    .vert0_valid_o         (valid_63_to_73_v0),
    .vert0_ready_i         (ready_73_to_63_v0),
    .vert1_data_i          (data_53_to_63_v1),
    .vert1_valid_i         (valid_53_to_63_v1),
    .vert1_ready_o         (ready_63_to_53_v1),
    .vert1_data_o          (data_63_to_73_v1),
    .vert1_valid_o         (valid_63_to_73_v1),
    .vert1_ready_i         (ready_73_to_63_v1),
    .local_data_i          (data_i[3][6]),
    .local_valid_i         (valid_i[3][6]),
    .local_ready_o         (ready_o[3][6]),
    .local_data_o          (data_o[3][6]),
    .local_valid_o         (valid_o[3][6]),
    .local_ready_i         (ready_i[3][6]),
    .credit_upd            (credit_upd)
);

/*Router 3,7*/    
cast_router #(
    .isUBM_list            (isUBM_list_3_7),
    .isFC_list             (isFC_list_3_7),
    .FCdn_list             (FCdn_list_3_7),
    .FCpl_list             (FCpl_list_3_7),
    .rt_file_list          (cast_rt_file_list_3_7)
)router_3_7(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_72_to_73),
    .west_valid_i          (valid_72_to_73),
    .west_ready_o          (ready_73_to_72),
    .west_data_o           (data_73_to_72),
    .west_valid_o          (valid_73_to_72),
    .west_ready_i          (ready_72_to_73),
    .east_data_i           (data_74_to_73),
    .east_valid_i          (valid_74_to_73),
    .east_ready_o          (ready_73_to_74),
    .east_data_o           (data_73_to_74),
    .east_valid_o          (valid_73_to_74),
    .east_ready_i          (ready_74_to_73),
    .vert0_data_i          (data_63_to_73_v0),
    .vert0_valid_i         (valid_63_to_73_v0),
    .vert0_ready_o         (ready_73_to_63_v0),
    .vert0_data_o          (data_73_to_83_v0),
    .vert0_valid_o         (valid_73_to_83_v0),
    .vert0_ready_i         (ready_83_to_73_v0),
    .vert1_data_i          (data_63_to_73_v1),
    .vert1_valid_i         (valid_63_to_73_v1),
    .vert1_ready_o         (ready_73_to_63_v1),
    .vert1_data_o          (data_73_to_83_v1),
    .vert1_valid_o         (valid_73_to_83_v1),
    .vert1_ready_i         (ready_83_to_73_v1),
    .local_data_i          (data_i[3][7]),
    .local_valid_i         (valid_i[3][7]),
    .local_ready_o         (ready_o[3][7]),
    .local_data_o          (data_o[3][7]),
    .local_valid_o         (valid_o[3][7]),
    .local_ready_i         (ready_i[3][7]),
    .credit_upd            (credit_upd)
);

/*Router 3,8*/    
cast_router #(
    .isUBM_list            (isUBM_list_3_8),
    .isFC_list             (isFC_list_3_8),
    .FCdn_list             (FCdn_list_3_8),
    .FCpl_list             (FCpl_list_3_8),
    .rt_file_list          (cast_rt_file_list_3_8)
)router_3_8(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_82_to_83),
    .west_valid_i          (valid_82_to_83),
    .west_ready_o          (ready_83_to_82),
    .west_data_o           (data_83_to_82),
    .west_valid_o          (valid_83_to_82),
    .west_ready_i          (ready_82_to_83),
    .east_data_i           (data_84_to_83),
    .east_valid_i          (valid_84_to_83),
    .east_ready_o          (ready_83_to_84),
    .east_data_o           (data_83_to_84),
    .east_valid_o          (valid_83_to_84),
    .east_ready_i          (ready_84_to_83),
    .vert0_data_i          (data_73_to_83_v0),
    .vert0_valid_i         (valid_73_to_83_v0),
    .vert0_ready_o         (ready_83_to_73_v0),
    .vert0_data_o          (data_83_to_93_v0),
    .vert0_valid_o         (valid_83_to_93_v0),
    .vert0_ready_i         (ready_93_to_83_v0),
    .vert1_data_i          (data_73_to_83_v1),
    .vert1_valid_i         (valid_73_to_83_v1),
    .vert1_ready_o         (ready_83_to_73_v1),
    .vert1_data_o          (data_83_to_93_v1),
    .vert1_valid_o         (valid_83_to_93_v1),
    .vert1_ready_i         (ready_93_to_83_v1),
    .local_data_i          (data_i[3][8]),
    .local_valid_i         (valid_i[3][8]),
    .local_ready_o         (ready_o[3][8]),
    .local_data_o          (data_o[3][8]),
    .local_valid_o         (valid_o[3][8]),
    .local_ready_i         (ready_i[3][8]),
    .credit_upd            (credit_upd)
);

/*Router 3,9*/    
cast_router #(
    .isUBM_list            (isUBM_list_3_9),
    .isFC_list             (isFC_list_3_9),
    .FCdn_list             (FCdn_list_3_9),
    .FCpl_list             (FCpl_list_3_9),
    .rt_file_list          (cast_rt_file_list_3_9)
)router_3_9(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_92_to_93),
    .west_valid_i          (valid_92_to_93),
    .west_ready_o          (ready_93_to_92),
    .west_data_o           (data_93_to_92),
    .west_valid_o          (valid_93_to_92),
    .west_ready_i          (ready_92_to_93),
    .east_data_i           (data_94_to_93),
    .east_valid_i          (valid_94_to_93),
    .east_ready_o          (ready_93_to_94),
    .east_data_o           (data_93_to_94),
    .east_valid_o          (valid_93_to_94),
    .east_ready_i          (ready_94_to_93),
    .vert0_data_i          (data_83_to_93_v0),
    .vert0_valid_i         (valid_83_to_93_v0),
    .vert0_ready_o         (ready_93_to_83_v0),
    .vert0_data_o          (data_93_to_103_v0),
    .vert0_valid_o         (valid_93_to_103_v0),
    .vert0_ready_i         (ready_103_to_93_v0),
    .vert1_data_i          (data_83_to_93_v1),
    .vert1_valid_i         (valid_83_to_93_v1),
    .vert1_ready_o         (ready_93_to_83_v1),
    .vert1_data_o          (data_93_to_103_v1),
    .vert1_valid_o         (valid_93_to_103_v1),
    .vert1_ready_i         (ready_103_to_93_v1),
    .local_data_i          (data_i[3][9]),
    .local_valid_i         (valid_i[3][9]),
    .local_ready_o         (ready_o[3][9]),
    .local_data_o          (data_o[3][9]),
    .local_valid_o         (valid_o[3][9]),
    .local_ready_i         (ready_i[3][9]),
    .credit_upd            (credit_upd)
);

/*Router 3,10*/    
cast_router #(
    .isUBM_list            (isUBM_list_3_10),
    .isFC_list             (isFC_list_3_10),
    .FCdn_list             (FCdn_list_3_10),
    .FCpl_list             (FCpl_list_3_10),
    .rt_file_list          (cast_rt_file_list_3_10)
)router_3_10(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_102_to_103),
    .west_valid_i          (valid_102_to_103),
    .west_ready_o          (ready_103_to_102),
    .west_data_o           (data_103_to_102),
    .west_valid_o          (valid_103_to_102),
    .west_ready_i          (ready_102_to_103),
    .east_data_i           (data_104_to_103),
    .east_valid_i          (valid_104_to_103),
    .east_ready_o          (ready_103_to_104),
    .east_data_o           (data_103_to_104),
    .east_valid_o          (valid_103_to_104),
    .east_ready_i          (ready_104_to_103),
    .vert0_data_i          (data_93_to_103_v0),
    .vert0_valid_i         (valid_93_to_103_v0),
    .vert0_ready_o         (ready_103_to_93_v0),
    .vert0_data_o          (data_103_to_113_v0),
    .vert0_valid_o         (valid_103_to_113_v0),
    .vert0_ready_i         (ready_113_to_103_v0),
    .vert1_data_i          (data_93_to_103_v1),
    .vert1_valid_i         (valid_93_to_103_v1),
    .vert1_ready_o         (ready_103_to_93_v1),
    .vert1_data_o          (data_103_to_113_v1),
    .vert1_valid_o         (valid_103_to_113_v1),
    .vert1_ready_i         (ready_113_to_103_v1),
    .local_data_i          (data_i[3][10]),
    .local_valid_i         (valid_i[3][10]),
    .local_ready_o         (ready_o[3][10]),
    .local_data_o          (data_o[3][10]),
    .local_valid_o         (valid_o[3][10]),
    .local_ready_i         (ready_i[3][10]),
    .credit_upd            (credit_upd)
);

/*Router 3,11*/    
cast_router #(
    .isUBM_list            (isUBM_list_3_11),
    .isFC_list             (isFC_list_3_11),
    .FCdn_list             (FCdn_list_3_11),
    .FCpl_list             (FCpl_list_3_11),
    .rt_file_list          (cast_rt_file_list_3_11)
)router_3_11(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_112_to_113),
    .west_valid_i          (valid_112_to_113),
    .west_ready_o          (ready_113_to_112),
    .west_data_o           (data_113_to_112),
    .west_valid_o          (valid_113_to_112),
    .west_ready_i          (ready_112_to_113),
    .east_data_i           (data_114_to_113),
    .east_valid_i          (valid_114_to_113),
    .east_ready_o          (ready_113_to_114),
    .east_data_o           (data_113_to_114),
    .east_valid_o          (valid_113_to_114),
    .east_ready_i          (ready_114_to_113),
    .vert0_data_i          (data_103_to_113_v0),
    .vert0_valid_i         (valid_103_to_113_v0),
    .vert0_ready_o         (ready_113_to_103_v0),
    .vert0_data_o          (data_113_to_123_v0),
    .vert0_valid_o         (valid_113_to_123_v0),
    .vert0_ready_i         (ready_123_to_113_v0),
    .vert1_data_i          (data_103_to_113_v1),
    .vert1_valid_i         (valid_103_to_113_v1),
    .vert1_ready_o         (ready_113_to_103_v1),
    .vert1_data_o          (data_113_to_123_v1),
    .vert1_valid_o         (valid_113_to_123_v1),
    .vert1_ready_i         (ready_123_to_113_v1),
    .local_data_i          (data_i[3][11]),
    .local_valid_i         (valid_i[3][11]),
    .local_ready_o         (ready_o[3][11]),
    .local_data_o          (data_o[3][11]),
    .local_valid_o         (valid_o[3][11]),
    .local_ready_i         (ready_i[3][11]),
    .credit_upd            (credit_upd)
);

/*Router 3,12*/    
cast_router #(
    .isUBM_list            (isUBM_list_3_12),
    .isFC_list             (isFC_list_3_12),
    .FCdn_list             (FCdn_list_3_12),
    .FCpl_list             (FCpl_list_3_12),
    .rt_file_list          (cast_rt_file_list_3_12)
)router_3_12(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_122_to_123),
    .west_valid_i          (valid_122_to_123),
    .west_ready_o          (ready_123_to_122),
    .west_data_o           (data_123_to_122),
    .west_valid_o          (valid_123_to_122),
    .west_ready_i          (ready_122_to_123),
    .east_data_i           (data_124_to_123),
    .east_valid_i          (valid_124_to_123),
    .east_ready_o          (ready_123_to_124),
    .east_data_o           (data_123_to_124),
    .east_valid_o          (valid_123_to_124),
    .east_ready_i          (ready_124_to_123),
    .vert0_data_i          (data_113_to_123_v0),
    .vert0_valid_i         (valid_113_to_123_v0),
    .vert0_ready_o         (ready_123_to_113_v0),
    .vert0_data_o          (data_123_to_133_v0),
    .vert0_valid_o         (valid_123_to_133_v0),
    .vert0_ready_i         (ready_133_to_123_v0),
    .vert1_data_i          (data_113_to_123_v1),
    .vert1_valid_i         (valid_113_to_123_v1),
    .vert1_ready_o         (ready_123_to_113_v1),
    .vert1_data_o          (data_123_to_133_v1),
    .vert1_valid_o         (valid_123_to_133_v1),
    .vert1_ready_i         (ready_133_to_123_v1),
    .local_data_i          (data_i[3][12]),
    .local_valid_i         (valid_i[3][12]),
    .local_ready_o         (ready_o[3][12]),
    .local_data_o          (data_o[3][12]),
    .local_valid_o         (valid_o[3][12]),
    .local_ready_i         (ready_i[3][12]),
    .credit_upd            (credit_upd)
);

/*Router 3,13*/    
cast_router #(
    .isUBM_list            (isUBM_list_3_13),
    .isFC_list             (isFC_list_3_13),
    .FCdn_list             (FCdn_list_3_13),
    .FCpl_list             (FCpl_list_3_13),
    .rt_file_list          (cast_rt_file_list_3_13)
)router_3_13(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_132_to_133),
    .west_valid_i          (valid_132_to_133),
    .west_ready_o          (ready_133_to_132),
    .west_data_o           (data_133_to_132),
    .west_valid_o          (valid_133_to_132),
    .west_ready_i          (ready_132_to_133),
    .east_data_i           (data_134_to_133),
    .east_valid_i          (valid_134_to_133),
    .east_ready_o          (ready_133_to_134),
    .east_data_o           (data_133_to_134),
    .east_valid_o          (valid_133_to_134),
    .east_ready_i          (ready_134_to_133),
    .vert0_data_i          (data_123_to_133_v0),
    .vert0_valid_i         (valid_123_to_133_v0),
    .vert0_ready_o         (ready_133_to_123_v0),
    .vert0_data_o          (data_133_to_143_v0),
    .vert0_valid_o         (valid_133_to_143_v0),
    .vert0_ready_i         (ready_143_to_133_v0),
    .vert1_data_i          (data_123_to_133_v1),
    .vert1_valid_i         (valid_123_to_133_v1),
    .vert1_ready_o         (ready_133_to_123_v1),
    .vert1_data_o          (data_133_to_143_v1),
    .vert1_valid_o         (valid_133_to_143_v1),
    .vert1_ready_i         (ready_143_to_133_v1),
    .local_data_i          (data_i[3][13]),
    .local_valid_i         (valid_i[3][13]),
    .local_ready_o         (ready_o[3][13]),
    .local_data_o          (data_o[3][13]),
    .local_valid_o         (valid_o[3][13]),
    .local_ready_i         (ready_i[3][13]),
    .credit_upd            (credit_upd)
);

/*Router 3,14*/    
cast_router #(
    .isUBM_list            (isUBM_list_3_14),
    .isFC_list             (isFC_list_3_14),
    .FCdn_list             (FCdn_list_3_14),
    .FCpl_list             (FCpl_list_3_14),
    .rt_file_list          (cast_rt_file_list_3_14)
)router_3_14(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_142_to_143),
    .west_valid_i          (valid_142_to_143),
    .west_ready_o          (ready_143_to_142),
    .west_data_o           (data_143_to_142),
    .west_valid_o          (valid_143_to_142),
    .west_ready_i          (ready_142_to_143),
    .east_data_i           (data_144_to_143),
    .east_valid_i          (valid_144_to_143),
    .east_ready_o          (ready_143_to_144),
    .east_data_o           (data_143_to_144),
    .east_valid_o          (valid_143_to_144),
    .east_ready_i          (ready_144_to_143),
    .vert0_data_i          (data_133_to_143_v0),
    .vert0_valid_i         (valid_133_to_143_v0),
    .vert0_ready_o         (ready_143_to_133_v0),
    .vert0_data_o          (data_143_to_153_v0),
    .vert0_valid_o         (valid_143_to_153_v0),
    .vert0_ready_i         (ready_153_to_143_v0),
    .vert1_data_i          (data_133_to_143_v1),
    .vert1_valid_i         (valid_133_to_143_v1),
    .vert1_ready_o         (ready_143_to_133_v1),
    .vert1_data_o          (data_143_to_153_v1),
    .vert1_valid_o         (valid_143_to_153_v1),
    .vert1_ready_i         (ready_153_to_143_v1),
    .local_data_i          (data_i[3][14]),
    .local_valid_i         (valid_i[3][14]),
    .local_ready_o         (ready_o[3][14]),
    .local_data_o          (data_o[3][14]),
    .local_valid_o         (valid_o[3][14]),
    .local_ready_i         (ready_i[3][14]),
    .credit_upd            (credit_upd)
);

/*Router 3,15*/    
cast_router #(
    .isUBM_list            (isUBM_list_3_15),
    .isFC_list             (isFC_list_3_15),
    .FCdn_list             (FCdn_list_3_15),
    .FCpl_list             (FCpl_list_3_15),
    .rt_file_list          (cast_rt_file_list_3_15)
)router_3_15(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_152_to_153),
    .west_valid_i          (valid_152_to_153),
    .west_ready_o          (ready_153_to_152),
    .west_data_o           (data_153_to_152),
    .west_valid_o          (valid_153_to_152),
    .west_ready_i          (ready_152_to_153),
    .east_data_i           (data_154_to_153),
    .east_valid_i          (valid_154_to_153),
    .east_ready_o          (ready_153_to_154),
    .east_data_o           (data_153_to_154),
    .east_valid_o          (valid_153_to_154),
    .east_ready_i          (ready_154_to_153),
    .vert0_data_i          (data_143_to_153_v0),
    .vert0_valid_i         (valid_143_to_153_v0),
    .vert0_ready_o         (ready_153_to_143_v0),
    .vert0_data_o          (data_153_to_163_v0),
    .vert0_valid_o         (valid_153_to_163_v0),
    .vert0_ready_i         (ready_163_to_153_v0),
    .vert1_data_i          (data_143_to_153_v1),
    .vert1_valid_i         (valid_143_to_153_v1),
    .vert1_ready_o         (ready_153_to_143_v1),
    .vert1_data_o          (data_153_to_163_v1),
    .vert1_valid_o         (valid_153_to_163_v1),
    .vert1_ready_i         (ready_163_to_153_v1),
    .local_data_i          (data_i[3][15]),
    .local_valid_i         (valid_i[3][15]),
    .local_ready_o         (ready_o[3][15]),
    .local_data_o          (data_o[3][15]),
    .local_valid_o         (valid_o[3][15]),
    .local_ready_i         (ready_i[3][15]),
    .credit_upd            (credit_upd)
);

/*Router 3,16*/    
cast_router #(
    .isUBM_list            (isUBM_list_3_16),
    .isFC_list             (isFC_list_3_16),
    .FCdn_list             (FCdn_list_3_16),
    .FCpl_list             (FCpl_list_3_16),
    .rt_file_list          (cast_rt_file_list_3_16)
)router_3_16(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_162_to_163),
    .west_valid_i          (valid_162_to_163),
    .west_ready_o          (ready_163_to_162),
    .west_data_o           (data_163_to_162),
    .west_valid_o          (valid_163_to_162),
    .west_ready_i          (ready_162_to_163),
    .east_data_i           (data_164_to_163),
    .east_valid_i          (valid_164_to_163),
    .east_ready_o          (ready_163_to_164),
    .east_data_o           (data_163_to_164),
    .east_valid_o          (valid_163_to_164),
    .east_ready_i          (ready_164_to_163),
    .vert0_data_i          (data_153_to_163_v0),
    .vert0_valid_i         (valid_153_to_163_v0),
    .vert0_ready_o         (ready_163_to_153_v0),
    .vert0_data_o          (data_163_to_173_v0),
    .vert0_valid_o         (valid_163_to_173_v0),
    .vert0_ready_i         (ready_173_to_163_v0),
    .vert1_data_i          (data_153_to_163_v1),
    .vert1_valid_i         (valid_153_to_163_v1),
    .vert1_ready_o         (ready_163_to_153_v1),
    .vert1_data_o          (data_163_to_173_v1),
    .vert1_valid_o         (valid_163_to_173_v1),
    .vert1_ready_i         (ready_173_to_163_v1),
    .local_data_i          (data_i[3][16]),
    .local_valid_i         (valid_i[3][16]),
    .local_ready_o         (ready_o[3][16]),
    .local_data_o          (data_o[3][16]),
    .local_valid_o         (valid_o[3][16]),
    .local_ready_i         (ready_i[3][16]),
    .credit_upd            (credit_upd)
);

/*Router 3,17*/    
cast_router #(
    .isUBM_list            (isUBM_list_3_17),
    .isFC_list             (isFC_list_3_17),
    .FCdn_list             (FCdn_list_3_17),
    .FCpl_list             (FCpl_list_3_17),
    .rt_file_list          (cast_rt_file_list_3_17)
)router_3_17(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_172_to_173),
    .west_valid_i          (valid_172_to_173),
    .west_ready_o          (ready_173_to_172),
    .west_data_o           (data_173_to_172),
    .west_valid_o          (valid_173_to_172),
    .west_ready_i          (ready_172_to_173),
    .east_data_i           (data_174_to_173),
    .east_valid_i          (valid_174_to_173),
    .east_ready_o          (ready_173_to_174),
    .east_data_o           (data_173_to_174),
    .east_valid_o          (valid_173_to_174),
    .east_ready_i          (ready_174_to_173),
    .vert0_data_i          (data_163_to_173_v0),
    .vert0_valid_i         (valid_163_to_173_v0),
    .vert0_ready_o         (ready_173_to_163_v0),
    .vert0_data_o          (data_173_to_183_v0),
    .vert0_valid_o         (valid_173_to_183_v0),
    .vert0_ready_i         (ready_183_to_173_v0),
    .vert1_data_i          (data_163_to_173_v1),
    .vert1_valid_i         (valid_163_to_173_v1),
    .vert1_ready_o         (ready_173_to_163_v1),
    .vert1_data_o          (data_173_to_183_v1),
    .vert1_valid_o         (valid_173_to_183_v1),
    .vert1_ready_i         (ready_183_to_173_v1),
    .local_data_i          (data_i[3][17]),
    .local_valid_i         (valid_i[3][17]),
    .local_ready_o         (ready_o[3][17]),
    .local_data_o          (data_o[3][17]),
    .local_valid_o         (valid_o[3][17]),
    .local_ready_i         (ready_i[3][17]),
    .credit_upd            (credit_upd)
);

/*Router 3,18*/    
cast_router #(
    .isUBM_list            (isUBM_list_3_18),
    .isFC_list             (isFC_list_3_18),
    .FCdn_list             (FCdn_list_3_18),
    .FCpl_list             (FCpl_list_3_18),
    .rt_file_list          (cast_rt_file_list_3_18)
)router_3_18(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_182_to_183),
    .west_valid_i          (valid_182_to_183),
    .west_ready_o          (ready_183_to_182),
    .west_data_o           (data_183_to_182),
    .west_valid_o          (valid_183_to_182),
    .west_ready_i          (ready_182_to_183),
    .east_data_i           (data_184_to_183),
    .east_valid_i          (valid_184_to_183),
    .east_ready_o          (ready_183_to_184),
    .east_data_o           (data_183_to_184),
    .east_valid_o          (valid_183_to_184),
    .east_ready_i          (ready_184_to_183),
    .vert0_data_i          (data_173_to_183_v0),
    .vert0_valid_i         (valid_173_to_183_v0),
    .vert0_ready_o         (ready_183_to_173_v0),
    .vert0_data_o          (data_183_to_193_v0),
    .vert0_valid_o         (valid_183_to_193_v0),
    .vert0_ready_i         (ready_193_to_183_v0),
    .vert1_data_i          (data_173_to_183_v1),
    .vert1_valid_i         (valid_173_to_183_v1),
    .vert1_ready_o         (ready_183_to_173_v1),
    .vert1_data_o          (data_183_to_193_v1),
    .vert1_valid_o         (valid_183_to_193_v1),
    .vert1_ready_i         (ready_193_to_183_v1),
    .local_data_i          (data_i[3][18]),
    .local_valid_i         (valid_i[3][18]),
    .local_ready_o         (ready_o[3][18]),
    .local_data_o          (data_o[3][18]),
    .local_valid_o         (valid_o[3][18]),
    .local_ready_i         (ready_i[3][18]),
    .credit_upd            (credit_upd)
);

/*Router 3,19*/    
cast_router #(
    .isUBM_list            (isUBM_list_3_19),
    .isFC_list             (isFC_list_3_19),
    .FCdn_list             (FCdn_list_3_19),
    .FCpl_list             (FCpl_list_3_19),
    .rt_file_list          (cast_rt_file_list_3_19)
)router_3_19(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_192_to_193),
    .west_valid_i          (valid_192_to_193),
    .west_ready_o          (ready_193_to_192),
    .west_data_o           (data_193_to_192),
    .west_valid_o          (valid_193_to_192),
    .west_ready_i          (ready_192_to_193),
    .east_data_i           (data_194_to_193),
    .east_valid_i          (valid_194_to_193),
    .east_ready_o          (ready_193_to_194),
    .east_data_o           (data_193_to_194),
    .east_valid_o          (valid_193_to_194),
    .east_ready_i          (ready_194_to_193),
    .vert0_data_i          (data_183_to_193_v0),
    .vert0_valid_i         (valid_183_to_193_v0),
    .vert0_ready_o         (ready_193_to_183_v0),
    .vert0_data_o          (data_193_to_203_v0),
    .vert0_valid_o         (valid_193_to_203_v0),
    .vert0_ready_i         (ready_203_to_193_v0),
    .vert1_data_i          (data_183_to_193_v1),
    .vert1_valid_i         (valid_183_to_193_v1),
    .vert1_ready_o         (ready_193_to_183_v1),
    .vert1_data_o          (data_193_to_203_v1),
    .vert1_valid_o         (valid_193_to_203_v1),
    .vert1_ready_i         (ready_203_to_193_v1),
    .local_data_i          (data_i[3][19]),
    .local_valid_i         (valid_i[3][19]),
    .local_ready_o         (ready_o[3][19]),
    .local_data_o          (data_o[3][19]),
    .local_valid_o         (valid_o[3][19]),
    .local_ready_i         (ready_i[3][19]),
    .credit_upd            (credit_upd)
);

/*Router 3,20*/    
cast_router #(
    .isUBM_list            (isUBM_list_3_20),
    .isFC_list             (isFC_list_3_20),
    .FCdn_list             (FCdn_list_3_20),
    .FCpl_list             (FCpl_list_3_20),
    .rt_file_list          (cast_rt_file_list_3_20)
)router_3_20(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_202_to_203),
    .west_valid_i          (valid_202_to_203),
    .west_ready_o          (ready_203_to_202),
    .west_data_o           (data_203_to_202),
    .west_valid_o          (valid_203_to_202),
    .west_ready_i          (ready_202_to_203),
    .east_data_i           (data_204_to_203),
    .east_valid_i          (valid_204_to_203),
    .east_ready_o          (ready_203_to_204),
    .east_data_o           (data_203_to_204),
    .east_valid_o          (valid_203_to_204),
    .east_ready_i          (ready_204_to_203),
    .vert0_data_i          (data_193_to_203_v0),
    .vert0_valid_i         (valid_193_to_203_v0),
    .vert0_ready_o         (ready_203_to_193_v0),
    .vert0_data_o          (data_203_to_213_v0),
    .vert0_valid_o         (valid_203_to_213_v0),
    .vert0_ready_i         (ready_213_to_203_v0),
    .vert1_data_i          (data_193_to_203_v1),
    .vert1_valid_i         (valid_193_to_203_v1),
    .vert1_ready_o         (ready_203_to_193_v1),
    .vert1_data_o          (data_203_to_213_v1),
    .vert1_valid_o         (valid_203_to_213_v1),
    .vert1_ready_i         (ready_213_to_203_v1),
    .local_data_i          (data_i[3][20]),
    .local_valid_i         (valid_i[3][20]),
    .local_ready_o         (ready_o[3][20]),
    .local_data_o          (data_o[3][20]),
    .local_valid_o         (valid_o[3][20]),
    .local_ready_i         (ready_i[3][20]),
    .credit_upd            (credit_upd)
);

/*Router 3,21*/    
cast_router #(
    .isUBM_list            (isUBM_list_3_21),
    .isFC_list             (isFC_list_3_21),
    .FCdn_list             (FCdn_list_3_21),
    .FCpl_list             (FCpl_list_3_21),
    .rt_file_list          (cast_rt_file_list_3_21)
)router_3_21(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_212_to_213),
    .west_valid_i          (valid_212_to_213),
    .west_ready_o          (ready_213_to_212),
    .west_data_o           (data_213_to_212),
    .west_valid_o          (valid_213_to_212),
    .west_ready_i          (ready_212_to_213),
    .east_data_i           (data_214_to_213),
    .east_valid_i          (valid_214_to_213),
    .east_ready_o          (ready_213_to_214),
    .east_data_o           (data_213_to_214),
    .east_valid_o          (valid_213_to_214),
    .east_ready_i          (ready_214_to_213),
    .vert0_data_i          (data_203_to_213_v0),
    .vert0_valid_i         (valid_203_to_213_v0),
    .vert0_ready_o         (ready_213_to_203_v0),
    .vert0_data_o          (data_213_to_223_v0),
    .vert0_valid_o         (valid_213_to_223_v0),
    .vert0_ready_i         (ready_223_to_213_v0),
    .vert1_data_i          (data_203_to_213_v1),
    .vert1_valid_i         (valid_203_to_213_v1),
    .vert1_ready_o         (ready_213_to_203_v1),
    .vert1_data_o          (data_213_to_223_v1),
    .vert1_valid_o         (valid_213_to_223_v1),
    .vert1_ready_i         (ready_223_to_213_v1),
    .local_data_i          (data_i[3][21]),
    .local_valid_i         (valid_i[3][21]),
    .local_ready_o         (ready_o[3][21]),
    .local_data_o          (data_o[3][21]),
    .local_valid_o         (valid_o[3][21]),
    .local_ready_i         (ready_i[3][21]),
    .credit_upd            (credit_upd)
);

/*Router 3,22*/    
cast_router #(
    .isUBM_list            (isUBM_list_3_22),
    .isFC_list             (isFC_list_3_22),
    .FCdn_list             (FCdn_list_3_22),
    .FCpl_list             (FCpl_list_3_22),
    .rt_file_list          (cast_rt_file_list_3_22)
)router_3_22(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_222_to_223),
    .west_valid_i          (valid_222_to_223),
    .west_ready_o          (ready_223_to_222),
    .west_data_o           (data_223_to_222),
    .west_valid_o          (valid_223_to_222),
    .west_ready_i          (ready_222_to_223),
    .east_data_i           (data_224_to_223),
    .east_valid_i          (valid_224_to_223),
    .east_ready_o          (ready_223_to_224),
    .east_data_o           (data_223_to_224),
    .east_valid_o          (valid_223_to_224),
    .east_ready_i          (ready_224_to_223),
    .vert0_data_i          (data_213_to_223_v0),
    .vert0_valid_i         (valid_213_to_223_v0),
    .vert0_ready_o         (ready_223_to_213_v0),
    .vert0_data_o          (data_223_to_233_v0),
    .vert0_valid_o         (valid_223_to_233_v0),
    .vert0_ready_i         (ready_233_to_223_v0),
    .vert1_data_i          (data_213_to_223_v1),
    .vert1_valid_i         (valid_213_to_223_v1),
    .vert1_ready_o         (ready_223_to_213_v1),
    .vert1_data_o          (data_223_to_233_v1),
    .vert1_valid_o         (valid_223_to_233_v1),
    .vert1_ready_i         (ready_233_to_223_v1),
    .local_data_i          (data_i[3][22]),
    .local_valid_i         (valid_i[3][22]),
    .local_ready_o         (ready_o[3][22]),
    .local_data_o          (data_o[3][22]),
    .local_valid_o         (valid_o[3][22]),
    .local_ready_i         (ready_i[3][22]),
    .credit_upd            (credit_upd)
);

/*Router 3,23*/    
cast_router #(
    .isUBM_list            (isUBM_list_3_23),
    .isFC_list             (isFC_list_3_23),
    .FCdn_list             (FCdn_list_3_23),
    .FCpl_list             (FCpl_list_3_23),
    .rt_file_list          (cast_rt_file_list_3_23)
)router_3_23(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_232_to_233),
    .west_valid_i          (valid_232_to_233),
    .west_ready_o          (ready_233_to_232),
    .west_data_o           (data_o_flee5),
    .west_valid_o          (valid_o_flee5),
    .west_ready_i          (ready_i_flee5),
    .east_data_i           (data_234_to_233),
    .east_valid_i          (valid_234_to_233),
    .east_ready_o          (ready_233_to_234),
    .east_data_o           (data_233_to_234),
    .east_valid_o          (valid_233_to_234),
    .east_ready_i          (ready_234_to_233),
    .vert0_data_i          (data_223_to_233_v0),
    .vert0_valid_i         (valid_223_to_233_v0),
    .vert0_ready_o         (ready_233_to_223_v0),
    .vert0_data_o          (data_233_to_243_v0),
    .vert0_valid_o         (valid_233_to_243_v0),
    .vert0_ready_i         (ready_243_to_233_v0),
    .vert1_data_i          (data_223_to_233_v1),
    .vert1_valid_i         (valid_223_to_233_v1),
    .vert1_ready_o         (ready_233_to_223_v1),
    .vert1_data_o          (data_233_to_243_v1),
    .vert1_valid_o         (valid_233_to_243_v1),
    .vert1_ready_i         (ready_243_to_233_v1),
    .local_data_i          (data_i[3][23]),
    .local_valid_i         (valid_i[3][23]),
    .local_ready_o         (ready_o[3][23]),
    .local_data_o          (data_o[3][23]),
    .local_valid_o         (valid_o[3][23]),
    .local_ready_i         (ready_i[3][23]),
    .credit_upd            (credit_upd)
);

/*Router 3,24*/    
cast_router #(
    .isUBM_list            (isUBM_list_3_24),
    .isFC_list             (isFC_list_3_24),
    .FCdn_list             (FCdn_list_3_24),
    .FCpl_list             (FCpl_list_3_24),
    .rt_file_list          (cast_rt_file_list_3_24)
)router_3_24(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_242_to_243),
    .west_valid_i          (valid_242_to_243),
    .west_ready_o          (ready_243_to_242),
    .west_data_o           (data_243_to_242),
    .west_valid_o          (valid_243_to_242),
    .west_ready_i          (ready_242_to_243),
    .east_data_i           (data_244_to_243),
    .east_valid_i          (valid_244_to_243),
    .east_ready_o          (ready_243_to_244),
    .east_data_o           (data_243_to_244),
    .east_valid_o          (valid_243_to_244),
    .east_ready_i          (ready_244_to_243),
    .vert0_data_i          (data_233_to_243_v0),
    .vert0_valid_i         (valid_233_to_243_v0),
    .vert0_ready_o         (ready_243_to_233_v0),
    .vert0_data_o          (),
    .vert0_valid_o         (),
    .vert0_ready_i         (1'b0),
    .vert1_data_i          (data_233_to_243_v1),
    .vert1_valid_i         (valid_233_to_243_v1),
    .vert1_ready_o         (ready_243_to_233_v1),
    .vert1_data_o          (),
    .vert1_valid_o         (),
    .vert1_ready_i         (1'b0),
    .local_data_i          (data_i[3][24]),
    .local_valid_i         (valid_i[3][24]),
    .local_ready_o         (ready_o[3][24]),
    .local_data_o          (data_o[3][24]),
    .local_valid_o         (valid_o[3][24]),
    .local_ready_i         (ready_i[3][24]),
    .credit_upd            (credit_upd)
);

/*Router 4,0*/    
cast_router #(
    .isUBM_list            (isUBM_list_4_0),
    .isFC_list             (isFC_list_4_0),
    .FCdn_list             (FCdn_list_4_0),
    .FCpl_list             (FCpl_list_4_0),
    .rt_file_list          (cast_rt_file_list_4_0)
)router_4_0(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_3_to_4),
    .west_valid_i          (valid_3_to_4),
    .west_ready_o          (ready_4_to_3),
    .west_data_o           (data_4_to_3),
    .west_valid_o          (valid_4_to_3),
    .west_ready_i          (ready_3_to_4),
    .east_data_i           (data_5_to_4),
    .east_valid_i          (valid_5_to_4),
    .east_ready_o          (ready_4_to_5),
    .east_data_o           (data_4_to_5),
    .east_valid_o          (valid_4_to_5),
    .east_ready_i          (ready_5_to_4),
    .vert0_data_i          (34'b0),
    .vert0_valid_i         (1'b0),
    .vert0_ready_o         (),
    .vert0_data_o          (data_4_to_14_v0),
    .vert0_valid_o         (valid_4_to_14_v0),
    .vert0_ready_i         (ready_14_to_4_v0),
    .vert1_data_i          (34'b0),
    .vert1_valid_i         (1'b0),
    .vert1_ready_o         (),
    .vert1_data_o          (data_4_to_14_v1),
    .vert1_valid_o         (valid_4_to_14_v1),
    .vert1_ready_i         (ready_14_to_4_v1),
    .local_data_i          (data_i[4][0]),
    .local_valid_i         (valid_i[4][0]),
    .local_ready_o         (ready_o[4][0]),
    .local_data_o          (data_o[4][0]),
    .local_valid_o         (valid_o[4][0]),
    .local_ready_i         (ready_i[4][0]),
    .credit_upd            (credit_upd)
);

/*Router 4,1*/    
cast_router #(
    .isUBM_list            (isUBM_list_4_1),
    .isFC_list             (isFC_list_4_1),
    .FCdn_list             (FCdn_list_4_1),
    .FCpl_list             (FCpl_list_4_1),
    .rt_file_list          (cast_rt_file_list_4_1)
)router_4_1(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_13_to_14),
    .west_valid_i          (valid_13_to_14),
    .west_ready_o          (ready_14_to_13),
    .west_data_o           (data_14_to_13),
    .west_valid_o          (valid_14_to_13),
    .west_ready_i          (ready_13_to_14),
    .east_data_i           (data_15_to_14),
    .east_valid_i          (valid_15_to_14),
    .east_ready_o          (ready_14_to_15),
    .east_data_o           (data_14_to_15),
    .east_valid_o          (valid_14_to_15),
    .east_ready_i          (ready_15_to_14),
    .vert0_data_i          (data_4_to_14_v0),
    .vert0_valid_i         (valid_4_to_14_v0),
    .vert0_ready_o         (ready_14_to_4_v0),
    .vert0_data_o          (data_14_to_24_v0),
    .vert0_valid_o         (valid_14_to_24_v0),
    .vert0_ready_i         (ready_24_to_14_v0),
    .vert1_data_i          (data_4_to_14_v1),
    .vert1_valid_i         (valid_4_to_14_v1),
    .vert1_ready_o         (ready_14_to_4_v1),
    .vert1_data_o          (data_14_to_24_v1),
    .vert1_valid_o         (valid_14_to_24_v1),
    .vert1_ready_i         (ready_24_to_14_v1),
    .local_data_i          (data_i[4][1]),
    .local_valid_i         (valid_i[4][1]),
    .local_ready_o         (ready_o[4][1]),
    .local_data_o          (data_o[4][1]),
    .local_valid_o         (valid_o[4][1]),
    .local_ready_i         (ready_i[4][1]),
    .credit_upd            (credit_upd)
);

/*Router 4,2*/    
cast_router #(
    .isUBM_list            (isUBM_list_4_2),
    .isFC_list             (isFC_list_4_2),
    .FCdn_list             (FCdn_list_4_2),
    .FCpl_list             (FCpl_list_4_2),
    .rt_file_list          (cast_rt_file_list_4_2)
)router_4_2(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_23_to_24),
    .west_valid_i          (valid_23_to_24),
    .west_ready_o          (ready_24_to_23),
    .west_data_o           (data_24_to_23),
    .west_valid_o          (valid_24_to_23),
    .west_ready_i          (ready_23_to_24),
    .east_data_i           (data_25_to_24),
    .east_valid_i          (valid_25_to_24),
    .east_ready_o          (ready_24_to_25),
    .east_data_o           (data_24_to_25),
    .east_valid_o          (valid_24_to_25),
    .east_ready_i          (ready_25_to_24),
    .vert0_data_i          (data_14_to_24_v0),
    .vert0_valid_i         (valid_14_to_24_v0),
    .vert0_ready_o         (ready_24_to_14_v0),
    .vert0_data_o          (data_24_to_34_v0),
    .vert0_valid_o         (valid_24_to_34_v0),
    .vert0_ready_i         (ready_34_to_24_v0),
    .vert1_data_i          (data_14_to_24_v1),
    .vert1_valid_i         (valid_14_to_24_v1),
    .vert1_ready_o         (ready_24_to_14_v1),
    .vert1_data_o          (data_24_to_34_v1),
    .vert1_valid_o         (valid_24_to_34_v1),
    .vert1_ready_i         (ready_34_to_24_v1),
    .local_data_i          (data_i[4][2]),
    .local_valid_i         (valid_i[4][2]),
    .local_ready_o         (ready_o[4][2]),
    .local_data_o          (data_o[4][2]),
    .local_valid_o         (valid_o[4][2]),
    .local_ready_i         (ready_i[4][2]),
    .credit_upd            (credit_upd)
);

/*Router 4,3*/    
cast_router #(
    .isUBM_list            (isUBM_list_4_3),
    .isFC_list             (isFC_list_4_3),
    .FCdn_list             (FCdn_list_4_3),
    .FCpl_list             (FCpl_list_4_3),
    .rt_file_list          (cast_rt_file_list_4_3)
)router_4_3(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_33_to_34),
    .west_valid_i          (valid_33_to_34),
    .west_ready_o          (ready_34_to_33),
    .west_data_o           (data_34_to_33),
    .west_valid_o          (valid_34_to_33),
    .west_ready_i          (ready_33_to_34),
    .east_data_i           (data_35_to_34),
    .east_valid_i          (valid_35_to_34),
    .east_ready_o          (ready_34_to_35),
    .east_data_o           (data_34_to_35),
    .east_valid_o          (valid_34_to_35),
    .east_ready_i          (ready_35_to_34),
    .vert0_data_i          (data_24_to_34_v0),
    .vert0_valid_i         (valid_24_to_34_v0),
    .vert0_ready_o         (ready_34_to_24_v0),
    .vert0_data_o          (data_34_to_44_v0),
    .vert0_valid_o         (valid_34_to_44_v0),
    .vert0_ready_i         (ready_44_to_34_v0),
    .vert1_data_i          (data_24_to_34_v1),
    .vert1_valid_i         (valid_24_to_34_v1),
    .vert1_ready_o         (ready_34_to_24_v1),
    .vert1_data_o          (data_34_to_44_v1),
    .vert1_valid_o         (valid_34_to_44_v1),
    .vert1_ready_i         (ready_44_to_34_v1),
    .local_data_i          (data_i[4][3]),
    .local_valid_i         (valid_i[4][3]),
    .local_ready_o         (ready_o[4][3]),
    .local_data_o          (data_o[4][3]),
    .local_valid_o         (valid_o[4][3]),
    .local_ready_i         (ready_i[4][3]),
    .credit_upd            (credit_upd)
);

/*Router 4,4*/    
cast_router #(
    .isUBM_list            (isUBM_list_4_4),
    .isFC_list             (isFC_list_4_4),
    .FCdn_list             (FCdn_list_4_4),
    .FCpl_list             (FCpl_list_4_4),
    .rt_file_list          (cast_rt_file_list_4_4)
)router_4_4(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_43_to_44),
    .west_valid_i          (valid_43_to_44),
    .west_ready_o          (ready_44_to_43),
    .west_data_o           (data_44_to_43),
    .west_valid_o          (valid_44_to_43),
    .west_ready_i          (ready_43_to_44),
    .east_data_i           (data_45_to_44),
    .east_valid_i          (valid_45_to_44),
    .east_ready_o          (ready_44_to_45),
    .east_data_o           (data_44_to_45),
    .east_valid_o          (valid_44_to_45),
    .east_ready_i          (ready_45_to_44),
    .vert0_data_i          (data_34_to_44_v0),
    .vert0_valid_i         (valid_34_to_44_v0),
    .vert0_ready_o         (ready_44_to_34_v0),
    .vert0_data_o          (data_44_to_54_v0),
    .vert0_valid_o         (valid_44_to_54_v0),
    .vert0_ready_i         (ready_54_to_44_v0),
    .vert1_data_i          (data_34_to_44_v1),
    .vert1_valid_i         (valid_34_to_44_v1),
    .vert1_ready_o         (ready_44_to_34_v1),
    .vert1_data_o          (data_44_to_54_v1),
    .vert1_valid_o         (valid_44_to_54_v1),
    .vert1_ready_i         (ready_54_to_44_v1),
    .local_data_i          (data_i[4][4]),
    .local_valid_i         (valid_i[4][4]),
    .local_ready_o         (ready_o[4][4]),
    .local_data_o          (data_o[4][4]),
    .local_valid_o         (valid_o[4][4]),
    .local_ready_i         (ready_i[4][4]),
    .credit_upd            (credit_upd)
);

/*Router 4,5*/    
cast_router #(
    .isUBM_list            (isUBM_list_4_5),
    .isFC_list             (isFC_list_4_5),
    .FCdn_list             (FCdn_list_4_5),
    .FCpl_list             (FCpl_list_4_5),
    .rt_file_list          (cast_rt_file_list_4_5)
)router_4_5(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_53_to_54),
    .west_valid_i          (valid_53_to_54),
    .west_ready_o          (ready_54_to_53),
    .west_data_o           (data_54_to_53),
    .west_valid_o          (valid_54_to_53),
    .west_ready_i          (ready_53_to_54),
    .east_data_i           (data_55_to_54),
    .east_valid_i          (valid_55_to_54),
    .east_ready_o          (ready_54_to_55),
    .east_data_o           (data_54_to_55),
    .east_valid_o          (valid_54_to_55),
    .east_ready_i          (ready_55_to_54),
    .vert0_data_i          (data_44_to_54_v0),
    .vert0_valid_i         (valid_44_to_54_v0),
    .vert0_ready_o         (ready_54_to_44_v0),
    .vert0_data_o          (data_54_to_64_v0),
    .vert0_valid_o         (valid_54_to_64_v0),
    .vert0_ready_i         (ready_64_to_54_v0),
    .vert1_data_i          (data_44_to_54_v1),
    .vert1_valid_i         (valid_44_to_54_v1),
    .vert1_ready_o         (ready_54_to_44_v1),
    .vert1_data_o          (data_54_to_64_v1),
    .vert1_valid_o         (valid_54_to_64_v1),
    .vert1_ready_i         (ready_64_to_54_v1),
    .local_data_i          (data_i[4][5]),
    .local_valid_i         (valid_i[4][5]),
    .local_ready_o         (ready_o[4][5]),
    .local_data_o          (data_o[4][5]),
    .local_valid_o         (valid_o[4][5]),
    .local_ready_i         (ready_i[4][5]),
    .credit_upd            (credit_upd)
);

/*Router 4,6*/    
cast_router #(
    .isUBM_list            (isUBM_list_4_6),
    .isFC_list             (isFC_list_4_6),
    .FCdn_list             (FCdn_list_4_6),
    .FCpl_list             (FCpl_list_4_6),
    .rt_file_list          (cast_rt_file_list_4_6)
)router_4_6(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_63_to_64),
    .west_valid_i          (valid_63_to_64),
    .west_ready_o          (ready_64_to_63),
    .west_data_o           (data_64_to_63),
    .west_valid_o          (valid_64_to_63),
    .west_ready_i          (ready_63_to_64),
    .east_data_i           (data_65_to_64),
    .east_valid_i          (valid_65_to_64),
    .east_ready_o          (ready_64_to_65),
    .east_data_o           (data_64_to_65),
    .east_valid_o          (valid_64_to_65),
    .east_ready_i          (ready_65_to_64),
    .vert0_data_i          (data_54_to_64_v0),
    .vert0_valid_i         (valid_54_to_64_v0),
    .vert0_ready_o         (ready_64_to_54_v0),
    .vert0_data_o          (data_64_to_74_v0),
    .vert0_valid_o         (valid_64_to_74_v0),
    .vert0_ready_i         (ready_74_to_64_v0),
    .vert1_data_i          (data_54_to_64_v1),
    .vert1_valid_i         (valid_54_to_64_v1),
    .vert1_ready_o         (ready_64_to_54_v1),
    .vert1_data_o          (data_64_to_74_v1),
    .vert1_valid_o         (valid_64_to_74_v1),
    .vert1_ready_i         (ready_74_to_64_v1),
    .local_data_i          (data_i[4][6]),
    .local_valid_i         (valid_i[4][6]),
    .local_ready_o         (ready_o[4][6]),
    .local_data_o          (data_o[4][6]),
    .local_valid_o         (valid_o[4][6]),
    .local_ready_i         (ready_i[4][6]),
    .credit_upd            (credit_upd)
);

/*Router 4,7*/    
cast_router #(
    .isUBM_list            (isUBM_list_4_7),
    .isFC_list             (isFC_list_4_7),
    .FCdn_list             (FCdn_list_4_7),
    .FCpl_list             (FCpl_list_4_7),
    .rt_file_list          (cast_rt_file_list_4_7)
)router_4_7(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_73_to_74),
    .west_valid_i          (valid_73_to_74),
    .west_ready_o          (ready_74_to_73),
    .west_data_o           (data_74_to_73),
    .west_valid_o          (valid_74_to_73),
    .west_ready_i          (ready_73_to_74),
    .east_data_i           (data_75_to_74),
    .east_valid_i          (valid_75_to_74),
    .east_ready_o          (ready_74_to_75),
    .east_data_o           (data_74_to_75),
    .east_valid_o          (valid_74_to_75),
    .east_ready_i          (ready_75_to_74),
    .vert0_data_i          (data_64_to_74_v0),
    .vert0_valid_i         (valid_64_to_74_v0),
    .vert0_ready_o         (ready_74_to_64_v0),
    .vert0_data_o          (data_74_to_84_v0),
    .vert0_valid_o         (valid_74_to_84_v0),
    .vert0_ready_i         (ready_84_to_74_v0),
    .vert1_data_i          (data_64_to_74_v1),
    .vert1_valid_i         (valid_64_to_74_v1),
    .vert1_ready_o         (ready_74_to_64_v1),
    .vert1_data_o          (data_74_to_84_v1),
    .vert1_valid_o         (valid_74_to_84_v1),
    .vert1_ready_i         (ready_84_to_74_v1),
    .local_data_i          (data_i[4][7]),
    .local_valid_i         (valid_i[4][7]),
    .local_ready_o         (ready_o[4][7]),
    .local_data_o          (data_o[4][7]),
    .local_valid_o         (valid_o[4][7]),
    .local_ready_i         (ready_i[4][7]),
    .credit_upd            (credit_upd)
);

/*Router 4,8*/    
cast_router #(
    .isUBM_list            (isUBM_list_4_8),
    .isFC_list             (isFC_list_4_8),
    .FCdn_list             (FCdn_list_4_8),
    .FCpl_list             (FCpl_list_4_8),
    .rt_file_list          (cast_rt_file_list_4_8)
)router_4_8(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_83_to_84),
    .west_valid_i          (valid_83_to_84),
    .west_ready_o          (ready_84_to_83),
    .west_data_o           (data_84_to_83),
    .west_valid_o          (valid_84_to_83),
    .west_ready_i          (ready_83_to_84),
    .east_data_i           (data_85_to_84),
    .east_valid_i          (valid_85_to_84),
    .east_ready_o          (ready_84_to_85),
    .east_data_o           (data_84_to_85),
    .east_valid_o          (valid_84_to_85),
    .east_ready_i          (ready_85_to_84),
    .vert0_data_i          (data_74_to_84_v0),
    .vert0_valid_i         (valid_74_to_84_v0),
    .vert0_ready_o         (ready_84_to_74_v0),
    .vert0_data_o          (data_84_to_94_v0),
    .vert0_valid_o         (valid_84_to_94_v0),
    .vert0_ready_i         (ready_94_to_84_v0),
    .vert1_data_i          (data_74_to_84_v1),
    .vert1_valid_i         (valid_74_to_84_v1),
    .vert1_ready_o         (ready_84_to_74_v1),
    .vert1_data_o          (data_84_to_94_v1),
    .vert1_valid_o         (valid_84_to_94_v1),
    .vert1_ready_i         (ready_94_to_84_v1),
    .local_data_i          (data_i[4][8]),
    .local_valid_i         (valid_i[4][8]),
    .local_ready_o         (ready_o[4][8]),
    .local_data_o          (data_o[4][8]),
    .local_valid_o         (valid_o[4][8]),
    .local_ready_i         (ready_i[4][8]),
    .credit_upd            (credit_upd)
);

/*Router 4,9*/    
cast_router #(
    .isUBM_list            (isUBM_list_4_9),
    .isFC_list             (isFC_list_4_9),
    .FCdn_list             (FCdn_list_4_9),
    .FCpl_list             (FCpl_list_4_9),
    .rt_file_list          (cast_rt_file_list_4_9)
)router_4_9(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_93_to_94),
    .west_valid_i          (valid_93_to_94),
    .west_ready_o          (ready_94_to_93),
    .west_data_o           (data_94_to_93),
    .west_valid_o          (valid_94_to_93),
    .west_ready_i          (ready_93_to_94),
    .east_data_i           (data_95_to_94),
    .east_valid_i          (valid_95_to_94),
    .east_ready_o          (ready_94_to_95),
    .east_data_o           (data_94_to_95),
    .east_valid_o          (valid_94_to_95),
    .east_ready_i          (ready_95_to_94),
    .vert0_data_i          (data_84_to_94_v0),
    .vert0_valid_i         (valid_84_to_94_v0),
    .vert0_ready_o         (ready_94_to_84_v0),
    .vert0_data_o          (data_94_to_104_v0),
    .vert0_valid_o         (valid_94_to_104_v0),
    .vert0_ready_i         (ready_104_to_94_v0),
    .vert1_data_i          (data_84_to_94_v1),
    .vert1_valid_i         (valid_84_to_94_v1),
    .vert1_ready_o         (ready_94_to_84_v1),
    .vert1_data_o          (data_94_to_104_v1),
    .vert1_valid_o         (valid_94_to_104_v1),
    .vert1_ready_i         (ready_104_to_94_v1),
    .local_data_i          (data_i[4][9]),
    .local_valid_i         (valid_i[4][9]),
    .local_ready_o         (ready_o[4][9]),
    .local_data_o          (data_o[4][9]),
    .local_valid_o         (valid_o[4][9]),
    .local_ready_i         (ready_i[4][9]),
    .credit_upd            (credit_upd)
);

/*Router 4,10*/    
cast_router #(
    .isUBM_list            (isUBM_list_4_10),
    .isFC_list             (isFC_list_4_10),
    .FCdn_list             (FCdn_list_4_10),
    .FCpl_list             (FCpl_list_4_10),
    .rt_file_list          (cast_rt_file_list_4_10)
)router_4_10(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_103_to_104),
    .west_valid_i          (valid_103_to_104),
    .west_ready_o          (ready_104_to_103),
    .west_data_o           (data_104_to_103),
    .west_valid_o          (valid_104_to_103),
    .west_ready_i          (ready_103_to_104),
    .east_data_i           (data_105_to_104),
    .east_valid_i          (valid_105_to_104),
    .east_ready_o          (ready_104_to_105),
    .east_data_o           (data_104_to_105),
    .east_valid_o          (valid_104_to_105),
    .east_ready_i          (ready_105_to_104),
    .vert0_data_i          (data_94_to_104_v0),
    .vert0_valid_i         (valid_94_to_104_v0),
    .vert0_ready_o         (ready_104_to_94_v0),
    .vert0_data_o          (data_104_to_114_v0),
    .vert0_valid_o         (valid_104_to_114_v0),
    .vert0_ready_i         (ready_114_to_104_v0),
    .vert1_data_i          (data_94_to_104_v1),
    .vert1_valid_i         (valid_94_to_104_v1),
    .vert1_ready_o         (ready_104_to_94_v1),
    .vert1_data_o          (data_104_to_114_v1),
    .vert1_valid_o         (valid_104_to_114_v1),
    .vert1_ready_i         (ready_114_to_104_v1),
    .local_data_i          (data_i[4][10]),
    .local_valid_i         (valid_i[4][10]),
    .local_ready_o         (ready_o[4][10]),
    .local_data_o          (data_o[4][10]),
    .local_valid_o         (valid_o[4][10]),
    .local_ready_i         (ready_i[4][10]),
    .credit_upd            (credit_upd)
);

/*Router 4,11*/    
cast_router #(
    .isUBM_list            (isUBM_list_4_11),
    .isFC_list             (isFC_list_4_11),
    .FCdn_list             (FCdn_list_4_11),
    .FCpl_list             (FCpl_list_4_11),
    .rt_file_list          (cast_rt_file_list_4_11)
)router_4_11(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_113_to_114),
    .west_valid_i          (valid_113_to_114),
    .west_ready_o          (ready_114_to_113),
    .west_data_o           (data_114_to_113),
    .west_valid_o          (valid_114_to_113),
    .west_ready_i          (ready_113_to_114),
    .east_data_i           (data_115_to_114),
    .east_valid_i          (valid_115_to_114),
    .east_ready_o          (ready_114_to_115),
    .east_data_o           (data_114_to_115),
    .east_valid_o          (valid_114_to_115),
    .east_ready_i          (ready_115_to_114),
    .vert0_data_i          (data_104_to_114_v0),
    .vert0_valid_i         (valid_104_to_114_v0),
    .vert0_ready_o         (ready_114_to_104_v0),
    .vert0_data_o          (data_114_to_124_v0),
    .vert0_valid_o         (valid_114_to_124_v0),
    .vert0_ready_i         (ready_124_to_114_v0),
    .vert1_data_i          (data_104_to_114_v1),
    .vert1_valid_i         (valid_104_to_114_v1),
    .vert1_ready_o         (ready_114_to_104_v1),
    .vert1_data_o          (data_114_to_124_v1),
    .vert1_valid_o         (valid_114_to_124_v1),
    .vert1_ready_i         (ready_124_to_114_v1),
    .local_data_i          (data_i[4][11]),
    .local_valid_i         (valid_i[4][11]),
    .local_ready_o         (ready_o[4][11]),
    .local_data_o          (data_o[4][11]),
    .local_valid_o         (valid_o[4][11]),
    .local_ready_i         (ready_i[4][11]),
    .credit_upd            (credit_upd)
);

/*Router 4,12*/    
cast_router #(
    .isUBM_list            (isUBM_list_4_12),
    .isFC_list             (isFC_list_4_12),
    .FCdn_list             (FCdn_list_4_12),
    .FCpl_list             (FCpl_list_4_12),
    .rt_file_list          (cast_rt_file_list_4_12)
)router_4_12(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_123_to_124),
    .west_valid_i          (valid_123_to_124),
    .west_ready_o          (ready_124_to_123),
    .west_data_o           (data_124_to_123),
    .west_valid_o          (valid_124_to_123),
    .west_ready_i          (ready_123_to_124),
    .east_data_i           (data_125_to_124),
    .east_valid_i          (valid_125_to_124),
    .east_ready_o          (ready_124_to_125),
    .east_data_o           (data_124_to_125),
    .east_valid_o          (valid_124_to_125),
    .east_ready_i          (ready_125_to_124),
    .vert0_data_i          (data_114_to_124_v0),
    .vert0_valid_i         (valid_114_to_124_v0),
    .vert0_ready_o         (ready_124_to_114_v0),
    .vert0_data_o          (data_124_to_134_v0),
    .vert0_valid_o         (valid_124_to_134_v0),
    .vert0_ready_i         (ready_134_to_124_v0),
    .vert1_data_i          (data_114_to_124_v1),
    .vert1_valid_i         (valid_114_to_124_v1),
    .vert1_ready_o         (ready_124_to_114_v1),
    .vert1_data_o          (data_124_to_134_v1),
    .vert1_valid_o         (valid_124_to_134_v1),
    .vert1_ready_i         (ready_134_to_124_v1),
    .local_data_i          (data_i[4][12]),
    .local_valid_i         (valid_i[4][12]),
    .local_ready_o         (ready_o[4][12]),
    .local_data_o          (data_o[4][12]),
    .local_valid_o         (valid_o[4][12]),
    .local_ready_i         (ready_i[4][12]),
    .credit_upd            (credit_upd)
);

/*Router 4,13*/    
cast_router #(
    .isUBM_list            (isUBM_list_4_13),
    .isFC_list             (isFC_list_4_13),
    .FCdn_list             (FCdn_list_4_13),
    .FCpl_list             (FCpl_list_4_13),
    .rt_file_list          (cast_rt_file_list_4_13)
)router_4_13(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_133_to_134),
    .west_valid_i          (valid_133_to_134),
    .west_ready_o          (ready_134_to_133),
    .west_data_o           (data_134_to_133),
    .west_valid_o          (valid_134_to_133),
    .west_ready_i          (ready_133_to_134),
    .east_data_i           (data_135_to_134),
    .east_valid_i          (valid_135_to_134),
    .east_ready_o          (ready_134_to_135),
    .east_data_o           (data_134_to_135),
    .east_valid_o          (valid_134_to_135),
    .east_ready_i          (ready_135_to_134),
    .vert0_data_i          (data_124_to_134_v0),
    .vert0_valid_i         (valid_124_to_134_v0),
    .vert0_ready_o         (ready_134_to_124_v0),
    .vert0_data_o          (data_134_to_144_v0),
    .vert0_valid_o         (valid_134_to_144_v0),
    .vert0_ready_i         (ready_144_to_134_v0),
    .vert1_data_i          (data_124_to_134_v1),
    .vert1_valid_i         (valid_124_to_134_v1),
    .vert1_ready_o         (ready_134_to_124_v1),
    .vert1_data_o          (data_134_to_144_v1),
    .vert1_valid_o         (valid_134_to_144_v1),
    .vert1_ready_i         (ready_144_to_134_v1),
    .local_data_i          (data_i[4][13]),
    .local_valid_i         (valid_i[4][13]),
    .local_ready_o         (ready_o[4][13]),
    .local_data_o          (data_o[4][13]),
    .local_valid_o         (valid_o[4][13]),
    .local_ready_i         (ready_i[4][13]),
    .credit_upd            (credit_upd)
);

/*Router 4,14*/    
cast_router #(
    .isUBM_list            (isUBM_list_4_14),
    .isFC_list             (isFC_list_4_14),
    .FCdn_list             (FCdn_list_4_14),
    .FCpl_list             (FCpl_list_4_14),
    .rt_file_list          (cast_rt_file_list_4_14)
)router_4_14(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_143_to_144),
    .west_valid_i          (valid_143_to_144),
    .west_ready_o          (ready_144_to_143),
    .west_data_o           (data_144_to_143),
    .west_valid_o          (valid_144_to_143),
    .west_ready_i          (ready_143_to_144),
    .east_data_i           (data_145_to_144),
    .east_valid_i          (valid_145_to_144),
    .east_ready_o          (ready_144_to_145),
    .east_data_o           (data_144_to_145),
    .east_valid_o          (valid_144_to_145),
    .east_ready_i          (ready_145_to_144),
    .vert0_data_i          (data_134_to_144_v0),
    .vert0_valid_i         (valid_134_to_144_v0),
    .vert0_ready_o         (ready_144_to_134_v0),
    .vert0_data_o          (data_144_to_154_v0),
    .vert0_valid_o         (valid_144_to_154_v0),
    .vert0_ready_i         (ready_154_to_144_v0),
    .vert1_data_i          (data_134_to_144_v1),
    .vert1_valid_i         (valid_134_to_144_v1),
    .vert1_ready_o         (ready_144_to_134_v1),
    .vert1_data_o          (data_144_to_154_v1),
    .vert1_valid_o         (valid_144_to_154_v1),
    .vert1_ready_i         (ready_154_to_144_v1),
    .local_data_i          (data_i[4][14]),
    .local_valid_i         (valid_i[4][14]),
    .local_ready_o         (ready_o[4][14]),
    .local_data_o          (data_o[4][14]),
    .local_valid_o         (valid_o[4][14]),
    .local_ready_i         (ready_i[4][14]),
    .credit_upd            (credit_upd)
);

/*Router 4,15*/    
cast_router #(
    .isUBM_list            (isUBM_list_4_15),
    .isFC_list             (isFC_list_4_15),
    .FCdn_list             (FCdn_list_4_15),
    .FCpl_list             (FCpl_list_4_15),
    .rt_file_list          (cast_rt_file_list_4_15)
)router_4_15(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_153_to_154),
    .west_valid_i          (valid_153_to_154),
    .west_ready_o          (ready_154_to_153),
    .west_data_o           (data_154_to_153),
    .west_valid_o          (valid_154_to_153),
    .west_ready_i          (ready_153_to_154),
    .east_data_i           (data_155_to_154),
    .east_valid_i          (valid_155_to_154),
    .east_ready_o          (ready_154_to_155),
    .east_data_o           (data_154_to_155),
    .east_valid_o          (valid_154_to_155),
    .east_ready_i          (ready_155_to_154),
    .vert0_data_i          (data_144_to_154_v0),
    .vert0_valid_i         (valid_144_to_154_v0),
    .vert0_ready_o         (ready_154_to_144_v0),
    .vert0_data_o          (data_154_to_164_v0),
    .vert0_valid_o         (valid_154_to_164_v0),
    .vert0_ready_i         (ready_164_to_154_v0),
    .vert1_data_i          (data_144_to_154_v1),
    .vert1_valid_i         (valid_144_to_154_v1),
    .vert1_ready_o         (ready_154_to_144_v1),
    .vert1_data_o          (data_154_to_164_v1),
    .vert1_valid_o         (valid_154_to_164_v1),
    .vert1_ready_i         (ready_164_to_154_v1),
    .local_data_i          (data_i[4][15]),
    .local_valid_i         (valid_i[4][15]),
    .local_ready_o         (ready_o[4][15]),
    .local_data_o          (data_o[4][15]),
    .local_valid_o         (valid_o[4][15]),
    .local_ready_i         (ready_i[4][15]),
    .credit_upd            (credit_upd)
);

/*Router 4,16*/    
cast_router #(
    .isUBM_list            (isUBM_list_4_16),
    .isFC_list             (isFC_list_4_16),
    .FCdn_list             (FCdn_list_4_16),
    .FCpl_list             (FCpl_list_4_16),
    .rt_file_list          (cast_rt_file_list_4_16)
)router_4_16(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_163_to_164),
    .west_valid_i          (valid_163_to_164),
    .west_ready_o          (ready_164_to_163),
    .west_data_o           (data_164_to_163),
    .west_valid_o          (valid_164_to_163),
    .west_ready_i          (ready_163_to_164),
    .east_data_i           (data_165_to_164),
    .east_valid_i          (valid_165_to_164),
    .east_ready_o          (ready_164_to_165),
    .east_data_o           (data_164_to_165),
    .east_valid_o          (valid_164_to_165),
    .east_ready_i          (ready_165_to_164),
    .vert0_data_i          (data_154_to_164_v0),
    .vert0_valid_i         (valid_154_to_164_v0),
    .vert0_ready_o         (ready_164_to_154_v0),
    .vert0_data_o          (data_164_to_174_v0),
    .vert0_valid_o         (valid_164_to_174_v0),
    .vert0_ready_i         (ready_174_to_164_v0),
    .vert1_data_i          (data_154_to_164_v1),
    .vert1_valid_i         (valid_154_to_164_v1),
    .vert1_ready_o         (ready_164_to_154_v1),
    .vert1_data_o          (data_164_to_174_v1),
    .vert1_valid_o         (valid_164_to_174_v1),
    .vert1_ready_i         (ready_174_to_164_v1),
    .local_data_i          (data_i[4][16]),
    .local_valid_i         (valid_i[4][16]),
    .local_ready_o         (ready_o[4][16]),
    .local_data_o          (data_o[4][16]),
    .local_valid_o         (valid_o[4][16]),
    .local_ready_i         (ready_i[4][16]),
    .credit_upd            (credit_upd)
);

/*Router 4,17*/    
cast_router #(
    .isUBM_list            (isUBM_list_4_17),
    .isFC_list             (isFC_list_4_17),
    .FCdn_list             (FCdn_list_4_17),
    .FCpl_list             (FCpl_list_4_17),
    .rt_file_list          (cast_rt_file_list_4_17)
)router_4_17(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_173_to_174),
    .west_valid_i          (valid_173_to_174),
    .west_ready_o          (ready_174_to_173),
    .west_data_o           (data_174_to_173),
    .west_valid_o          (valid_174_to_173),
    .west_ready_i          (ready_173_to_174),
    .east_data_i           (data_175_to_174),
    .east_valid_i          (valid_175_to_174),
    .east_ready_o          (ready_174_to_175),
    .east_data_o           (data_174_to_175),
    .east_valid_o          (valid_174_to_175),
    .east_ready_i          (ready_175_to_174),
    .vert0_data_i          (data_164_to_174_v0),
    .vert0_valid_i         (valid_164_to_174_v0),
    .vert0_ready_o         (ready_174_to_164_v0),
    .vert0_data_o          (data_174_to_184_v0),
    .vert0_valid_o         (valid_174_to_184_v0),
    .vert0_ready_i         (ready_184_to_174_v0),
    .vert1_data_i          (data_164_to_174_v1),
    .vert1_valid_i         (valid_164_to_174_v1),
    .vert1_ready_o         (ready_174_to_164_v1),
    .vert1_data_o          (data_174_to_184_v1),
    .vert1_valid_o         (valid_174_to_184_v1),
    .vert1_ready_i         (ready_184_to_174_v1),
    .local_data_i          (data_i[4][17]),
    .local_valid_i         (valid_i[4][17]),
    .local_ready_o         (ready_o[4][17]),
    .local_data_o          (data_o[4][17]),
    .local_valid_o         (valid_o[4][17]),
    .local_ready_i         (ready_i[4][17]),
    .credit_upd            (credit_upd)
);

/*Router 4,18*/    
cast_router #(
    .isUBM_list            (isUBM_list_4_18),
    .isFC_list             (isFC_list_4_18),
    .FCdn_list             (FCdn_list_4_18),
    .FCpl_list             (FCpl_list_4_18),
    .rt_file_list          (cast_rt_file_list_4_18)
)router_4_18(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_183_to_184),
    .west_valid_i          (valid_183_to_184),
    .west_ready_o          (ready_184_to_183),
    .west_data_o           (data_184_to_183),
    .west_valid_o          (valid_184_to_183),
    .west_ready_i          (ready_183_to_184),
    .east_data_i           (data_185_to_184),
    .east_valid_i          (valid_185_to_184),
    .east_ready_o          (ready_184_to_185),
    .east_data_o           (data_184_to_185),
    .east_valid_o          (valid_184_to_185),
    .east_ready_i          (ready_185_to_184),
    .vert0_data_i          (data_174_to_184_v0),
    .vert0_valid_i         (valid_174_to_184_v0),
    .vert0_ready_o         (ready_184_to_174_v0),
    .vert0_data_o          (data_184_to_194_v0),
    .vert0_valid_o         (valid_184_to_194_v0),
    .vert0_ready_i         (ready_194_to_184_v0),
    .vert1_data_i          (data_174_to_184_v1),
    .vert1_valid_i         (valid_174_to_184_v1),
    .vert1_ready_o         (ready_184_to_174_v1),
    .vert1_data_o          (data_184_to_194_v1),
    .vert1_valid_o         (valid_184_to_194_v1),
    .vert1_ready_i         (ready_194_to_184_v1),
    .local_data_i          (data_i[4][18]),
    .local_valid_i         (valid_i[4][18]),
    .local_ready_o         (ready_o[4][18]),
    .local_data_o          (data_o[4][18]),
    .local_valid_o         (valid_o[4][18]),
    .local_ready_i         (ready_i[4][18]),
    .credit_upd            (credit_upd)
);

/*Router 4,19*/    
cast_router #(
    .isUBM_list            (isUBM_list_4_19),
    .isFC_list             (isFC_list_4_19),
    .FCdn_list             (FCdn_list_4_19),
    .FCpl_list             (FCpl_list_4_19),
    .rt_file_list          (cast_rt_file_list_4_19)
)router_4_19(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_193_to_194),
    .west_valid_i          (valid_193_to_194),
    .west_ready_o          (ready_194_to_193),
    .west_data_o           (data_194_to_193),
    .west_valid_o          (valid_194_to_193),
    .west_ready_i          (ready_193_to_194),
    .east_data_i           (data_195_to_194),
    .east_valid_i          (valid_195_to_194),
    .east_ready_o          (ready_194_to_195),
    .east_data_o           (data_194_to_195),
    .east_valid_o          (valid_194_to_195),
    .east_ready_i          (ready_195_to_194),
    .vert0_data_i          (data_184_to_194_v0),
    .vert0_valid_i         (valid_184_to_194_v0),
    .vert0_ready_o         (ready_194_to_184_v0),
    .vert0_data_o          (data_194_to_204_v0),
    .vert0_valid_o         (valid_194_to_204_v0),
    .vert0_ready_i         (ready_204_to_194_v0),
    .vert1_data_i          (data_184_to_194_v1),
    .vert1_valid_i         (valid_184_to_194_v1),
    .vert1_ready_o         (ready_194_to_184_v1),
    .vert1_data_o          (data_194_to_204_v1),
    .vert1_valid_o         (valid_194_to_204_v1),
    .vert1_ready_i         (ready_204_to_194_v1),
    .local_data_i          (data_i[4][19]),
    .local_valid_i         (valid_i[4][19]),
    .local_ready_o         (ready_o[4][19]),
    .local_data_o          (data_o[4][19]),
    .local_valid_o         (valid_o[4][19]),
    .local_ready_i         (ready_i[4][19]),
    .credit_upd            (credit_upd)
);

/*Router 4,20*/    
cast_router #(
    .isUBM_list            (isUBM_list_4_20),
    .isFC_list             (isFC_list_4_20),
    .FCdn_list             (FCdn_list_4_20),
    .FCpl_list             (FCpl_list_4_20),
    .rt_file_list          (cast_rt_file_list_4_20)
)router_4_20(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_203_to_204),
    .west_valid_i          (valid_203_to_204),
    .west_ready_o          (ready_204_to_203),
    .west_data_o           (data_204_to_203),
    .west_valid_o          (valid_204_to_203),
    .west_ready_i          (ready_203_to_204),
    .east_data_i           (data_205_to_204),
    .east_valid_i          (valid_205_to_204),
    .east_ready_o          (ready_204_to_205),
    .east_data_o           (data_204_to_205),
    .east_valid_o          (valid_204_to_205),
    .east_ready_i          (ready_205_to_204),
    .vert0_data_i          (data_194_to_204_v0),
    .vert0_valid_i         (valid_194_to_204_v0),
    .vert0_ready_o         (ready_204_to_194_v0),
    .vert0_data_o          (data_204_to_214_v0),
    .vert0_valid_o         (valid_204_to_214_v0),
    .vert0_ready_i         (ready_214_to_204_v0),
    .vert1_data_i          (data_194_to_204_v1),
    .vert1_valid_i         (valid_194_to_204_v1),
    .vert1_ready_o         (ready_204_to_194_v1),
    .vert1_data_o          (data_204_to_214_v1),
    .vert1_valid_o         (valid_204_to_214_v1),
    .vert1_ready_i         (ready_214_to_204_v1),
    .local_data_i          (data_i[4][20]),
    .local_valid_i         (valid_i[4][20]),
    .local_ready_o         (ready_o[4][20]),
    .local_data_o          (data_o[4][20]),
    .local_valid_o         (valid_o[4][20]),
    .local_ready_i         (ready_i[4][20]),
    .credit_upd            (credit_upd)
);

/*Router 4,21*/    
cast_router #(
    .isUBM_list            (isUBM_list_4_21),
    .isFC_list             (isFC_list_4_21),
    .FCdn_list             (FCdn_list_4_21),
    .FCpl_list             (FCpl_list_4_21),
    .rt_file_list          (cast_rt_file_list_4_21)
)router_4_21(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_213_to_214),
    .west_valid_i          (valid_213_to_214),
    .west_ready_o          (ready_214_to_213),
    .west_data_o           (data_214_to_213),
    .west_valid_o          (valid_214_to_213),
    .west_ready_i          (ready_213_to_214),
    .east_data_i           (data_215_to_214),
    .east_valid_i          (valid_215_to_214),
    .east_ready_o          (ready_214_to_215),
    .east_data_o           (data_214_to_215),
    .east_valid_o          (valid_214_to_215),
    .east_ready_i          (ready_215_to_214),
    .vert0_data_i          (data_204_to_214_v0),
    .vert0_valid_i         (valid_204_to_214_v0),
    .vert0_ready_o         (ready_214_to_204_v0),
    .vert0_data_o          (data_214_to_224_v0),
    .vert0_valid_o         (valid_214_to_224_v0),
    .vert0_ready_i         (ready_224_to_214_v0),
    .vert1_data_i          (data_204_to_214_v1),
    .vert1_valid_i         (valid_204_to_214_v1),
    .vert1_ready_o         (ready_214_to_204_v1),
    .vert1_data_o          (data_214_to_224_v1),
    .vert1_valid_o         (valid_214_to_224_v1),
    .vert1_ready_i         (ready_224_to_214_v1),
    .local_data_i          (data_i[4][21]),
    .local_valid_i         (valid_i[4][21]),
    .local_ready_o         (ready_o[4][21]),
    .local_data_o          (data_o[4][21]),
    .local_valid_o         (valid_o[4][21]),
    .local_ready_i         (ready_i[4][21]),
    .credit_upd            (credit_upd)
);

/*Router 4,22*/    
cast_router #(
    .isUBM_list            (isUBM_list_4_22),
    .isFC_list             (isFC_list_4_22),
    .FCdn_list             (FCdn_list_4_22),
    .FCpl_list             (FCpl_list_4_22),
    .rt_file_list          (cast_rt_file_list_4_22)
)router_4_22(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_223_to_224),
    .west_valid_i          (valid_223_to_224),
    .west_ready_o          (ready_224_to_223),
    .west_data_o           (data_224_to_223),
    .west_valid_o          (valid_224_to_223),
    .west_ready_i          (ready_223_to_224),
    .east_data_i           (data_225_to_224),
    .east_valid_i          (valid_225_to_224),
    .east_ready_o          (ready_224_to_225),
    .east_data_o           (data_224_to_225),
    .east_valid_o          (valid_224_to_225),
    .east_ready_i          (ready_225_to_224),
    .vert0_data_i          (data_214_to_224_v0),
    .vert0_valid_i         (valid_214_to_224_v0),
    .vert0_ready_o         (ready_224_to_214_v0),
    .vert0_data_o          (data_224_to_234_v0),
    .vert0_valid_o         (valid_224_to_234_v0),
    .vert0_ready_i         (ready_234_to_224_v0),
    .vert1_data_i          (data_214_to_224_v1),
    .vert1_valid_i         (valid_214_to_224_v1),
    .vert1_ready_o         (ready_224_to_214_v1),
    .vert1_data_o          (data_224_to_234_v1),
    .vert1_valid_o         (valid_224_to_234_v1),
    .vert1_ready_i         (ready_234_to_224_v1),
    .local_data_i          (data_i[4][22]),
    .local_valid_i         (valid_i[4][22]),
    .local_ready_o         (ready_o[4][22]),
    .local_data_o          (data_o[4][22]),
    .local_valid_o         (valid_o[4][22]),
    .local_ready_i         (ready_i[4][22]),
    .credit_upd            (credit_upd)
);

/*Router 4,23*/    
cast_router #(
    .isUBM_list            (isUBM_list_4_23),
    .isFC_list             (isFC_list_4_23),
    .FCdn_list             (FCdn_list_4_23),
    .FCpl_list             (FCpl_list_4_23),
    .rt_file_list          (cast_rt_file_list_4_23)
)router_4_23(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_233_to_234),
    .west_valid_i          (valid_233_to_234),
    .west_ready_o          (ready_234_to_233),
    .west_data_o           (data_234_to_233),
    .west_valid_o          (valid_234_to_233),
    .west_ready_i          (ready_233_to_234),
    .east_data_i           (data_235_to_234),
    .east_valid_i          (valid_235_to_234),
    .east_ready_o          (ready_234_to_235),
    .east_data_o           (data_234_to_235),
    .east_valid_o          (valid_234_to_235),
    .east_ready_i          (ready_235_to_234),
    .vert0_data_i          (data_224_to_234_v0),
    .vert0_valid_i         (valid_224_to_234_v0),
    .vert0_ready_o         (ready_234_to_224_v0),
    .vert0_data_o          (data_234_to_244_v0),
    .vert0_valid_o         (valid_234_to_244_v0),
    .vert0_ready_i         (ready_244_to_234_v0),
    .vert1_data_i          (data_224_to_234_v1),
    .vert1_valid_i         (valid_224_to_234_v1),
    .vert1_ready_o         (ready_234_to_224_v1),
    .vert1_data_o          (data_234_to_244_v1),
    .vert1_valid_o         (valid_234_to_244_v1),
    .vert1_ready_i         (ready_244_to_234_v1),
    .local_data_i          (data_i[4][23]),
    .local_valid_i         (valid_i[4][23]),
    .local_ready_o         (ready_o[4][23]),
    .local_data_o          (data_o[4][23]),
    .local_valid_o         (valid_o[4][23]),
    .local_ready_i         (ready_i[4][23]),
    .credit_upd            (credit_upd)
);

/*Router 4,24*/    
cast_router #(
    .isUBM_list            (isUBM_list_4_24),
    .isFC_list             (isFC_list_4_24),
    .FCdn_list             (FCdn_list_4_24),
    .FCpl_list             (FCpl_list_4_24),
    .rt_file_list          (cast_rt_file_list_4_24)
)router_4_24(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_243_to_244),
    .west_valid_i          (valid_243_to_244),
    .west_ready_o          (ready_244_to_243),
    .west_data_o           (data_244_to_243),
    .west_valid_o          (valid_244_to_243),
    .west_ready_i          (ready_243_to_244),
    .east_data_i           (data_245_to_244),
    .east_valid_i          (valid_245_to_244),
    .east_ready_o          (ready_244_to_245),
    .east_data_o           (data_244_to_245),
    .east_valid_o          (valid_244_to_245),
    .east_ready_i          (ready_245_to_244),
    .vert0_data_i          (data_234_to_244_v0),
    .vert0_valid_i         (valid_234_to_244_v0),
    .vert0_ready_o         (ready_244_to_234_v0),
    .vert0_data_o          (),
    .vert0_valid_o         (),
    .vert0_ready_i         (1'b0),
    .vert1_data_i          (data_234_to_244_v1),
    .vert1_valid_i         (valid_234_to_244_v1),
    .vert1_ready_o         (ready_244_to_234_v1),
    .vert1_data_o          (),
    .vert1_valid_o         (),
    .vert1_ready_i         (1'b0),
    .local_data_i          (data_i[4][24]),
    .local_valid_i         (valid_i[4][24]),
    .local_ready_o         (ready_o[4][24]),
    .local_data_o          (data_o[4][24]),
    .local_valid_o         (valid_o[4][24]),
    .local_ready_i         (ready_i[4][24]),
    .credit_upd            (credit_upd)
);

/*Router 5,0*/    
cast_router #(
    .isUBM_list            (isUBM_list_5_0),
    .isFC_list             (isFC_list_5_0),
    .FCdn_list             (FCdn_list_5_0),
    .FCpl_list             (FCpl_list_5_0),
    .rt_file_list          (cast_rt_file_list_5_0)
)router_5_0(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_4_to_5),
    .west_valid_i          (valid_4_to_5),
    .west_ready_o          (ready_5_to_4),
    .west_data_o           (data_5_to_4),
    .west_valid_o          (valid_5_to_4),
    .west_ready_i          (ready_4_to_5),
    .east_data_i           (data_6_to_5),
    .east_valid_i          (valid_6_to_5),
    .east_ready_o          (ready_5_to_6),
    .east_data_o           (data_5_to_6),
    .east_valid_o          (valid_5_to_6),
    .east_ready_i          (ready_6_to_5),
    .vert0_data_i          (34'b0),
    .vert0_valid_i         (1'b0),
    .vert0_ready_o         (),
    .vert0_data_o          (data_5_to_15_v0),
    .vert0_valid_o         (valid_5_to_15_v0),
    .vert0_ready_i         (ready_15_to_5_v0),
    .vert1_data_i          (34'b0),
    .vert1_valid_i         (1'b0),
    .vert1_ready_o         (),
    .vert1_data_o          (data_5_to_15_v1),
    .vert1_valid_o         (valid_5_to_15_v1),
    .vert1_ready_i         (ready_15_to_5_v1),
    .local_data_i          (data_i[5][0]),
    .local_valid_i         (valid_i[5][0]),
    .local_ready_o         (ready_o[5][0]),
    .local_data_o          (data_o[5][0]),
    .local_valid_o         (valid_o[5][0]),
    .local_ready_i         (ready_i[5][0]),
    .credit_upd            (credit_upd)
);

/*Router 5,1*/    
cast_router #(
    .isUBM_list            (isUBM_list_5_1),
    .isFC_list             (isFC_list_5_1),
    .FCdn_list             (FCdn_list_5_1),
    .FCpl_list             (FCpl_list_5_1),
    .rt_file_list          (cast_rt_file_list_5_1)
)router_5_1(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_14_to_15),
    .west_valid_i          (valid_14_to_15),
    .west_ready_o          (ready_15_to_14),
    .west_data_o           (data_15_to_14),
    .west_valid_o          (valid_15_to_14),
    .west_ready_i          (ready_14_to_15),
    .east_data_i           (data_16_to_15),
    .east_valid_i          (valid_16_to_15),
    .east_ready_o          (ready_15_to_16),
    .east_data_o           (data_15_to_16),
    .east_valid_o          (valid_15_to_16),
    .east_ready_i          (ready_16_to_15),
    .vert0_data_i          (data_5_to_15_v0),
    .vert0_valid_i         (valid_5_to_15_v0),
    .vert0_ready_o         (ready_15_to_5_v0),
    .vert0_data_o          (data_15_to_25_v0),
    .vert0_valid_o         (valid_15_to_25_v0),
    .vert0_ready_i         (ready_25_to_15_v0),
    .vert1_data_i          (data_5_to_15_v1),
    .vert1_valid_i         (valid_5_to_15_v1),
    .vert1_ready_o         (ready_15_to_5_v1),
    .vert1_data_o          (data_15_to_25_v1),
    .vert1_valid_o         (valid_15_to_25_v1),
    .vert1_ready_i         (ready_25_to_15_v1),
    .local_data_i          (data_i[5][1]),
    .local_valid_i         (valid_i[5][1]),
    .local_ready_o         (ready_o[5][1]),
    .local_data_o          (data_o[5][1]),
    .local_valid_o         (valid_o[5][1]),
    .local_ready_i         (ready_i[5][1]),
    .credit_upd            (credit_upd)
);

/*Router 5,2*/    
cast_router #(
    .isUBM_list            (isUBM_list_5_2),
    .isFC_list             (isFC_list_5_2),
    .FCdn_list             (FCdn_list_5_2),
    .FCpl_list             (FCpl_list_5_2),
    .rt_file_list          (cast_rt_file_list_5_2)
)router_5_2(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_24_to_25),
    .west_valid_i          (valid_24_to_25),
    .west_ready_o          (ready_25_to_24),
    .west_data_o           (data_25_to_24),
    .west_valid_o          (valid_25_to_24),
    .west_ready_i          (ready_24_to_25),
    .east_data_i           (data_26_to_25),
    .east_valid_i          (valid_26_to_25),
    .east_ready_o          (ready_25_to_26),
    .east_data_o           (data_25_to_26),
    .east_valid_o          (valid_25_to_26),
    .east_ready_i          (ready_26_to_25),
    .vert0_data_i          (data_15_to_25_v0),
    .vert0_valid_i         (valid_15_to_25_v0),
    .vert0_ready_o         (ready_25_to_15_v0),
    .vert0_data_o          (data_25_to_35_v0),
    .vert0_valid_o         (valid_25_to_35_v0),
    .vert0_ready_i         (ready_35_to_25_v0),
    .vert1_data_i          (data_15_to_25_v1),
    .vert1_valid_i         (valid_15_to_25_v1),
    .vert1_ready_o         (ready_25_to_15_v1),
    .vert1_data_o          (data_25_to_35_v1),
    .vert1_valid_o         (valid_25_to_35_v1),
    .vert1_ready_i         (ready_35_to_25_v1),
    .local_data_i          (data_i[5][2]),
    .local_valid_i         (valid_i[5][2]),
    .local_ready_o         (ready_o[5][2]),
    .local_data_o          (data_o[5][2]),
    .local_valid_o         (valid_o[5][2]),
    .local_ready_i         (ready_i[5][2]),
    .credit_upd            (credit_upd)
);

/*Router 5,3*/    
cast_router #(
    .isUBM_list            (isUBM_list_5_3),
    .isFC_list             (isFC_list_5_3),
    .FCdn_list             (FCdn_list_5_3),
    .FCpl_list             (FCpl_list_5_3),
    .rt_file_list          (cast_rt_file_list_5_3)
)router_5_3(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_34_to_35),
    .west_valid_i          (valid_34_to_35),
    .west_ready_o          (ready_35_to_34),
    .west_data_o           (data_35_to_34),
    .west_valid_o          (valid_35_to_34),
    .west_ready_i          (ready_34_to_35),
    .east_data_i           (data_36_to_35),
    .east_valid_i          (valid_36_to_35),
    .east_ready_o          (ready_35_to_36),
    .east_data_o           (data_35_to_36),
    .east_valid_o          (valid_35_to_36),
    .east_ready_i          (ready_36_to_35),
    .vert0_data_i          (data_25_to_35_v0),
    .vert0_valid_i         (valid_25_to_35_v0),
    .vert0_ready_o         (ready_35_to_25_v0),
    .vert0_data_o          (data_35_to_45_v0),
    .vert0_valid_o         (valid_35_to_45_v0),
    .vert0_ready_i         (ready_45_to_35_v0),
    .vert1_data_i          (data_25_to_35_v1),
    .vert1_valid_i         (valid_25_to_35_v1),
    .vert1_ready_o         (ready_35_to_25_v1),
    .vert1_data_o          (data_35_to_45_v1),
    .vert1_valid_o         (valid_35_to_45_v1),
    .vert1_ready_i         (ready_45_to_35_v1),
    .local_data_i          (data_i[5][3]),
    .local_valid_i         (valid_i[5][3]),
    .local_ready_o         (ready_o[5][3]),
    .local_data_o          (data_o[5][3]),
    .local_valid_o         (valid_o[5][3]),
    .local_ready_i         (ready_i[5][3]),
    .credit_upd            (credit_upd)
);

/*Router 5,4*/    
cast_router #(
    .isUBM_list            (isUBM_list_5_4),
    .isFC_list             (isFC_list_5_4),
    .FCdn_list             (FCdn_list_5_4),
    .FCpl_list             (FCpl_list_5_4),
    .rt_file_list          (cast_rt_file_list_5_4)
)router_5_4(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_44_to_45),
    .west_valid_i          (valid_44_to_45),
    .west_ready_o          (ready_45_to_44),
    .west_data_o           (data_45_to_44),
    .west_valid_o          (valid_45_to_44),
    .west_ready_i          (ready_44_to_45),
    .east_data_i           (data_46_to_45),
    .east_valid_i          (valid_46_to_45),
    .east_ready_o          (ready_45_to_46),
    .east_data_o           (data_45_to_46),
    .east_valid_o          (valid_45_to_46),
    .east_ready_i          (ready_46_to_45),
    .vert0_data_i          (data_35_to_45_v0),
    .vert0_valid_i         (valid_35_to_45_v0),
    .vert0_ready_o         (ready_45_to_35_v0),
    .vert0_data_o          (data_45_to_55_v0),
    .vert0_valid_o         (valid_45_to_55_v0),
    .vert0_ready_i         (ready_55_to_45_v0),
    .vert1_data_i          (data_35_to_45_v1),
    .vert1_valid_i         (valid_35_to_45_v1),
    .vert1_ready_o         (ready_45_to_35_v1),
    .vert1_data_o          (data_45_to_55_v1),
    .vert1_valid_o         (valid_45_to_55_v1),
    .vert1_ready_i         (ready_55_to_45_v1),
    .local_data_i          (data_i[5][4]),
    .local_valid_i         (valid_i[5][4]),
    .local_ready_o         (ready_o[5][4]),
    .local_data_o          (data_o[5][4]),
    .local_valid_o         (valid_o[5][4]),
    .local_ready_i         (ready_i[5][4]),
    .credit_upd            (credit_upd)
);

/*Router 5,5*/    
cast_router #(
    .isUBM_list            (isUBM_list_5_5),
    .isFC_list             (isFC_list_5_5),
    .FCdn_list             (FCdn_list_5_5),
    .FCpl_list             (FCpl_list_5_5),
    .rt_file_list          (cast_rt_file_list_5_5)
)router_5_5(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_54_to_55),
    .west_valid_i          (valid_54_to_55),
    .west_ready_o          (ready_55_to_54),
    .west_data_o           (data_55_to_54),
    .west_valid_o          (valid_55_to_54),
    .west_ready_i          (ready_54_to_55),
    .east_data_i           (data_56_to_55),
    .east_valid_i          (valid_56_to_55),
    .east_ready_o          (ready_55_to_56),
    .east_data_o           (data_55_to_56),
    .east_valid_o          (valid_55_to_56),
    .east_ready_i          (ready_56_to_55),
    .vert0_data_i          (data_45_to_55_v0),
    .vert0_valid_i         (valid_45_to_55_v0),
    .vert0_ready_o         (ready_55_to_45_v0),
    .vert0_data_o          (data_55_to_65_v0),
    .vert0_valid_o         (valid_55_to_65_v0),
    .vert0_ready_i         (ready_65_to_55_v0),
    .vert1_data_i          (data_45_to_55_v1),
    .vert1_valid_i         (valid_45_to_55_v1),
    .vert1_ready_o         (ready_55_to_45_v1),
    .vert1_data_o          (data_55_to_65_v1),
    .vert1_valid_o         (valid_55_to_65_v1),
    .vert1_ready_i         (ready_65_to_55_v1),
    .local_data_i          (data_i[5][5]),
    .local_valid_i         (valid_i[5][5]),
    .local_ready_o         (ready_o[5][5]),
    .local_data_o          (data_o[5][5]),
    .local_valid_o         (valid_o[5][5]),
    .local_ready_i         (ready_i[5][5]),
    .credit_upd            (credit_upd)
);

/*Router 5,6*/    
cast_router #(
    .isUBM_list            (isUBM_list_5_6),
    .isFC_list             (isFC_list_5_6),
    .FCdn_list             (FCdn_list_5_6),
    .FCpl_list             (FCpl_list_5_6),
    .rt_file_list          (cast_rt_file_list_5_6)
)router_5_6(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_64_to_65),
    .west_valid_i          (valid_64_to_65),
    .west_ready_o          (ready_65_to_64),
    .west_data_o           (data_65_to_64),
    .west_valid_o          (valid_65_to_64),
    .west_ready_i          (ready_64_to_65),
    .east_data_i           (data_66_to_65),
    .east_valid_i          (valid_66_to_65),
    .east_ready_o          (ready_65_to_66),
    .east_data_o           (data_65_to_66),
    .east_valid_o          (valid_65_to_66),
    .east_ready_i          (ready_66_to_65),
    .vert0_data_i          (data_55_to_65_v0),
    .vert0_valid_i         (valid_55_to_65_v0),
    .vert0_ready_o         (ready_65_to_55_v0),
    .vert0_data_o          (data_65_to_75_v0),
    .vert0_valid_o         (valid_65_to_75_v0),
    .vert0_ready_i         (ready_75_to_65_v0),
    .vert1_data_i          (data_55_to_65_v1),
    .vert1_valid_i         (valid_55_to_65_v1),
    .vert1_ready_o         (ready_65_to_55_v1),
    .vert1_data_o          (data_65_to_75_v1),
    .vert1_valid_o         (valid_65_to_75_v1),
    .vert1_ready_i         (ready_75_to_65_v1),
    .local_data_i          (data_i[5][6]),
    .local_valid_i         (valid_i[5][6]),
    .local_ready_o         (ready_o[5][6]),
    .local_data_o          (data_o[5][6]),
    .local_valid_o         (valid_o[5][6]),
    .local_ready_i         (ready_i[5][6]),
    .credit_upd            (credit_upd)
);

/*Router 5,7*/    
cast_router #(
    .isUBM_list            (isUBM_list_5_7),
    .isFC_list             (isFC_list_5_7),
    .FCdn_list             (FCdn_list_5_7),
    .FCpl_list             (FCpl_list_5_7),
    .rt_file_list          (cast_rt_file_list_5_7)
)router_5_7(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_74_to_75),
    .west_valid_i          (valid_74_to_75),
    .west_ready_o          (ready_75_to_74),
    .west_data_o           (data_75_to_74),
    .west_valid_o          (valid_75_to_74),
    .west_ready_i          (ready_74_to_75),
    .east_data_i           (data_76_to_75),
    .east_valid_i          (valid_76_to_75),
    .east_ready_o          (ready_75_to_76),
    .east_data_o           (data_75_to_76),
    .east_valid_o          (valid_75_to_76),
    .east_ready_i          (ready_76_to_75),
    .vert0_data_i          (data_65_to_75_v0),
    .vert0_valid_i         (valid_65_to_75_v0),
    .vert0_ready_o         (ready_75_to_65_v0),
    .vert0_data_o          (data_75_to_85_v0),
    .vert0_valid_o         (valid_75_to_85_v0),
    .vert0_ready_i         (ready_85_to_75_v0),
    .vert1_data_i          (data_65_to_75_v1),
    .vert1_valid_i         (valid_65_to_75_v1),
    .vert1_ready_o         (ready_75_to_65_v1),
    .vert1_data_o          (data_75_to_85_v1),
    .vert1_valid_o         (valid_75_to_85_v1),
    .vert1_ready_i         (ready_85_to_75_v1),
    .local_data_i          (data_i[5][7]),
    .local_valid_i         (valid_i[5][7]),
    .local_ready_o         (ready_o[5][7]),
    .local_data_o          (data_o[5][7]),
    .local_valid_o         (valid_o[5][7]),
    .local_ready_i         (ready_i[5][7]),
    .credit_upd            (credit_upd)
);

/*Router 5,8*/    
cast_router #(
    .isUBM_list            (isUBM_list_5_8),
    .isFC_list             (isFC_list_5_8),
    .FCdn_list             (FCdn_list_5_8),
    .FCpl_list             (FCpl_list_5_8),
    .rt_file_list          (cast_rt_file_list_5_8)
)router_5_8(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_84_to_85),
    .west_valid_i          (valid_84_to_85),
    .west_ready_o          (ready_85_to_84),
    .west_data_o           (data_85_to_84),
    .west_valid_o          (valid_85_to_84),
    .west_ready_i          (ready_84_to_85),
    .east_data_i           (data_86_to_85),
    .east_valid_i          (valid_86_to_85),
    .east_ready_o          (ready_85_to_86),
    .east_data_o           (data_85_to_86),
    .east_valid_o          (valid_85_to_86),
    .east_ready_i          (ready_86_to_85),
    .vert0_data_i          (data_75_to_85_v0),
    .vert0_valid_i         (valid_75_to_85_v0),
    .vert0_ready_o         (ready_85_to_75_v0),
    .vert0_data_o          (data_85_to_95_v0),
    .vert0_valid_o         (valid_85_to_95_v0),
    .vert0_ready_i         (ready_95_to_85_v0),
    .vert1_data_i          (data_75_to_85_v1),
    .vert1_valid_i         (valid_75_to_85_v1),
    .vert1_ready_o         (ready_85_to_75_v1),
    .vert1_data_o          (data_85_to_95_v1),
    .vert1_valid_o         (valid_85_to_95_v1),
    .vert1_ready_i         (ready_95_to_85_v1),
    .local_data_i          (data_i[5][8]),
    .local_valid_i         (valid_i[5][8]),
    .local_ready_o         (ready_o[5][8]),
    .local_data_o          (data_o[5][8]),
    .local_valid_o         (valid_o[5][8]),
    .local_ready_i         (ready_i[5][8]),
    .credit_upd            (credit_upd)
);

/*Router 5,9*/    
cast_router #(
    .isUBM_list            (isUBM_list_5_9),
    .isFC_list             (isFC_list_5_9),
    .FCdn_list             (FCdn_list_5_9),
    .FCpl_list             (FCpl_list_5_9),
    .rt_file_list          (cast_rt_file_list_5_9)
)router_5_9(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_94_to_95),
    .west_valid_i          (valid_94_to_95),
    .west_ready_o          (ready_95_to_94),
    .west_data_o           (data_95_to_94),
    .west_valid_o          (valid_95_to_94),
    .west_ready_i          (ready_94_to_95),
    .east_data_i           (data_96_to_95),
    .east_valid_i          (valid_96_to_95),
    .east_ready_o          (ready_95_to_96),
    .east_data_o           (data_95_to_96),
    .east_valid_o          (valid_95_to_96),
    .east_ready_i          (ready_96_to_95),
    .vert0_data_i          (data_85_to_95_v0),
    .vert0_valid_i         (valid_85_to_95_v0),
    .vert0_ready_o         (ready_95_to_85_v0),
    .vert0_data_o          (data_95_to_105_v0),
    .vert0_valid_o         (valid_95_to_105_v0),
    .vert0_ready_i         (ready_105_to_95_v0),
    .vert1_data_i          (data_85_to_95_v1),
    .vert1_valid_i         (valid_85_to_95_v1),
    .vert1_ready_o         (ready_95_to_85_v1),
    .vert1_data_o          (data_95_to_105_v1),
    .vert1_valid_o         (valid_95_to_105_v1),
    .vert1_ready_i         (ready_105_to_95_v1),
    .local_data_i          (data_i[5][9]),
    .local_valid_i         (valid_i[5][9]),
    .local_ready_o         (ready_o[5][9]),
    .local_data_o          (data_o[5][9]),
    .local_valid_o         (valid_o[5][9]),
    .local_ready_i         (ready_i[5][9]),
    .credit_upd            (credit_upd)
);

/*Router 5,10*/    
cast_router #(
    .isUBM_list            (isUBM_list_5_10),
    .isFC_list             (isFC_list_5_10),
    .FCdn_list             (FCdn_list_5_10),
    .FCpl_list             (FCpl_list_5_10),
    .rt_file_list          (cast_rt_file_list_5_10)
)router_5_10(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_104_to_105),
    .west_valid_i          (valid_104_to_105),
    .west_ready_o          (ready_105_to_104),
    .west_data_o           (data_105_to_104),
    .west_valid_o          (valid_105_to_104),
    .west_ready_i          (ready_104_to_105),
    .east_data_i           (data_106_to_105),
    .east_valid_i          (valid_106_to_105),
    .east_ready_o          (ready_105_to_106),
    .east_data_o           (data_105_to_106),
    .east_valid_o          (valid_105_to_106),
    .east_ready_i          (ready_106_to_105),
    .vert0_data_i          (data_95_to_105_v0),
    .vert0_valid_i         (valid_95_to_105_v0),
    .vert0_ready_o         (ready_105_to_95_v0),
    .vert0_data_o          (data_105_to_115_v0),
    .vert0_valid_o         (valid_105_to_115_v0),
    .vert0_ready_i         (ready_115_to_105_v0),
    .vert1_data_i          (data_95_to_105_v1),
    .vert1_valid_i         (valid_95_to_105_v1),
    .vert1_ready_o         (ready_105_to_95_v1),
    .vert1_data_o          (data_105_to_115_v1),
    .vert1_valid_o         (valid_105_to_115_v1),
    .vert1_ready_i         (ready_115_to_105_v1),
    .local_data_i          (data_i[5][10]),
    .local_valid_i         (valid_i[5][10]),
    .local_ready_o         (ready_o[5][10]),
    .local_data_o          (data_o[5][10]),
    .local_valid_o         (valid_o[5][10]),
    .local_ready_i         (ready_i[5][10]),
    .credit_upd            (credit_upd)
);

/*Router 5,11*/    
cast_router #(
    .isUBM_list            (isUBM_list_5_11),
    .isFC_list             (isFC_list_5_11),
    .FCdn_list             (FCdn_list_5_11),
    .FCpl_list             (FCpl_list_5_11),
    .rt_file_list          (cast_rt_file_list_5_11)
)router_5_11(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_114_to_115),
    .west_valid_i          (valid_114_to_115),
    .west_ready_o          (ready_115_to_114),
    .west_data_o           (data_115_to_114),
    .west_valid_o          (valid_115_to_114),
    .west_ready_i          (ready_114_to_115),
    .east_data_i           (data_116_to_115),
    .east_valid_i          (valid_116_to_115),
    .east_ready_o          (ready_115_to_116),
    .east_data_o           (data_115_to_116),
    .east_valid_o          (valid_115_to_116),
    .east_ready_i          (ready_116_to_115),
    .vert0_data_i          (data_105_to_115_v0),
    .vert0_valid_i         (valid_105_to_115_v0),
    .vert0_ready_o         (ready_115_to_105_v0),
    .vert0_data_o          (data_115_to_125_v0),
    .vert0_valid_o         (valid_115_to_125_v0),
    .vert0_ready_i         (ready_125_to_115_v0),
    .vert1_data_i          (data_105_to_115_v1),
    .vert1_valid_i         (valid_105_to_115_v1),
    .vert1_ready_o         (ready_115_to_105_v1),
    .vert1_data_o          (data_115_to_125_v1),
    .vert1_valid_o         (valid_115_to_125_v1),
    .vert1_ready_i         (ready_125_to_115_v1),
    .local_data_i          (data_i[5][11]),
    .local_valid_i         (valid_i[5][11]),
    .local_ready_o         (ready_o[5][11]),
    .local_data_o          (data_o[5][11]),
    .local_valid_o         (valid_o[5][11]),
    .local_ready_i         (ready_i[5][11]),
    .credit_upd            (credit_upd)
);

/*Router 5,12*/    
cast_router #(
    .isUBM_list            (isUBM_list_5_12),
    .isFC_list             (isFC_list_5_12),
    .FCdn_list             (FCdn_list_5_12),
    .FCpl_list             (FCpl_list_5_12),
    .rt_file_list          (cast_rt_file_list_5_12)
)router_5_12(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_124_to_125),
    .west_valid_i          (valid_124_to_125),
    .west_ready_o          (ready_125_to_124),
    .west_data_o           (data_125_to_124),
    .west_valid_o          (valid_125_to_124),
    .west_ready_i          (ready_124_to_125),
    .east_data_i           (data_126_to_125),
    .east_valid_i          (valid_126_to_125),
    .east_ready_o          (ready_125_to_126),
    .east_data_o           (data_125_to_126),
    .east_valid_o          (valid_125_to_126),
    .east_ready_i          (ready_126_to_125),
    .vert0_data_i          (data_115_to_125_v0),
    .vert0_valid_i         (valid_115_to_125_v0),
    .vert0_ready_o         (ready_125_to_115_v0),
    .vert0_data_o          (data_125_to_135_v0),
    .vert0_valid_o         (valid_125_to_135_v0),
    .vert0_ready_i         (ready_135_to_125_v0),
    .vert1_data_i          (data_115_to_125_v1),
    .vert1_valid_i         (valid_115_to_125_v1),
    .vert1_ready_o         (ready_125_to_115_v1),
    .vert1_data_o          (data_125_to_135_v1),
    .vert1_valid_o         (valid_125_to_135_v1),
    .vert1_ready_i         (ready_135_to_125_v1),
    .local_data_i          (data_i[5][12]),
    .local_valid_i         (valid_i[5][12]),
    .local_ready_o         (ready_o[5][12]),
    .local_data_o          (data_o[5][12]),
    .local_valid_o         (valid_o[5][12]),
    .local_ready_i         (ready_i[5][12]),
    .credit_upd            (credit_upd)
);

/*Router 5,13*/    
cast_router #(
    .isUBM_list            (isUBM_list_5_13),
    .isFC_list             (isFC_list_5_13),
    .FCdn_list             (FCdn_list_5_13),
    .FCpl_list             (FCpl_list_5_13),
    .rt_file_list          (cast_rt_file_list_5_13)
)router_5_13(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_134_to_135),
    .west_valid_i          (valid_134_to_135),
    .west_ready_o          (ready_135_to_134),
    .west_data_o           (data_135_to_134),
    .west_valid_o          (valid_135_to_134),
    .west_ready_i          (ready_134_to_135),
    .east_data_i           (data_136_to_135),
    .east_valid_i          (valid_136_to_135),
    .east_ready_o          (ready_135_to_136),
    .east_data_o           (data_135_to_136),
    .east_valid_o          (valid_135_to_136),
    .east_ready_i          (ready_136_to_135),
    .vert0_data_i          (data_125_to_135_v0),
    .vert0_valid_i         (valid_125_to_135_v0),
    .vert0_ready_o         (ready_135_to_125_v0),
    .vert0_data_o          (data_135_to_145_v0),
    .vert0_valid_o         (valid_135_to_145_v0),
    .vert0_ready_i         (ready_145_to_135_v0),
    .vert1_data_i          (data_125_to_135_v1),
    .vert1_valid_i         (valid_125_to_135_v1),
    .vert1_ready_o         (ready_135_to_125_v1),
    .vert1_data_o          (data_135_to_145_v1),
    .vert1_valid_o         (valid_135_to_145_v1),
    .vert1_ready_i         (ready_145_to_135_v1),
    .local_data_i          (data_i[5][13]),
    .local_valid_i         (valid_i[5][13]),
    .local_ready_o         (ready_o[5][13]),
    .local_data_o          (data_o[5][13]),
    .local_valid_o         (valid_o[5][13]),
    .local_ready_i         (ready_i[5][13]),
    .credit_upd            (credit_upd)
);

/*Router 5,14*/    
cast_router #(
    .isUBM_list            (isUBM_list_5_14),
    .isFC_list             (isFC_list_5_14),
    .FCdn_list             (FCdn_list_5_14),
    .FCpl_list             (FCpl_list_5_14),
    .rt_file_list          (cast_rt_file_list_5_14)
)router_5_14(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_144_to_145),
    .west_valid_i          (valid_144_to_145),
    .west_ready_o          (ready_145_to_144),
    .west_data_o           (data_145_to_144),
    .west_valid_o          (valid_145_to_144),
    .west_ready_i          (ready_144_to_145),
    .east_data_i           (data_146_to_145),
    .east_valid_i          (valid_146_to_145),
    .east_ready_o          (ready_145_to_146),
    .east_data_o           (data_145_to_146),
    .east_valid_o          (valid_145_to_146),
    .east_ready_i          (ready_146_to_145),
    .vert0_data_i          (data_135_to_145_v0),
    .vert0_valid_i         (valid_135_to_145_v0),
    .vert0_ready_o         (ready_145_to_135_v0),
    .vert0_data_o          (data_145_to_155_v0),
    .vert0_valid_o         (valid_145_to_155_v0),
    .vert0_ready_i         (ready_155_to_145_v0),
    .vert1_data_i          (data_135_to_145_v1),
    .vert1_valid_i         (valid_135_to_145_v1),
    .vert1_ready_o         (ready_145_to_135_v1),
    .vert1_data_o          (data_145_to_155_v1),
    .vert1_valid_o         (valid_145_to_155_v1),
    .vert1_ready_i         (ready_155_to_145_v1),
    .local_data_i          (data_i[5][14]),
    .local_valid_i         (valid_i[5][14]),
    .local_ready_o         (ready_o[5][14]),
    .local_data_o          (data_o[5][14]),
    .local_valid_o         (valid_o[5][14]),
    .local_ready_i         (ready_i[5][14]),
    .credit_upd            (credit_upd)
);

/*Router 5,15*/    
cast_router #(
    .isUBM_list            (isUBM_list_5_15),
    .isFC_list             (isFC_list_5_15),
    .FCdn_list             (FCdn_list_5_15),
    .FCpl_list             (FCpl_list_5_15),
    .rt_file_list          (cast_rt_file_list_5_15)
)router_5_15(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_154_to_155),
    .west_valid_i          (valid_154_to_155),
    .west_ready_o          (ready_155_to_154),
    .west_data_o           (data_155_to_154),
    .west_valid_o          (valid_155_to_154),
    .west_ready_i          (ready_154_to_155),
    .east_data_i           (data_156_to_155),
    .east_valid_i          (valid_156_to_155),
    .east_ready_o          (ready_155_to_156),
    .east_data_o           (data_155_to_156),
    .east_valid_o          (valid_155_to_156),
    .east_ready_i          (ready_156_to_155),
    .vert0_data_i          (data_145_to_155_v0),
    .vert0_valid_i         (valid_145_to_155_v0),
    .vert0_ready_o         (ready_155_to_145_v0),
    .vert0_data_o          (data_155_to_165_v0),
    .vert0_valid_o         (valid_155_to_165_v0),
    .vert0_ready_i         (ready_165_to_155_v0),
    .vert1_data_i          (data_145_to_155_v1),
    .vert1_valid_i         (valid_145_to_155_v1),
    .vert1_ready_o         (ready_155_to_145_v1),
    .vert1_data_o          (data_155_to_165_v1),
    .vert1_valid_o         (valid_155_to_165_v1),
    .vert1_ready_i         (ready_165_to_155_v1),
    .local_data_i          (data_i[5][15]),
    .local_valid_i         (valid_i[5][15]),
    .local_ready_o         (ready_o[5][15]),
    .local_data_o          (data_o[5][15]),
    .local_valid_o         (valid_o[5][15]),
    .local_ready_i         (ready_i[5][15]),
    .credit_upd            (credit_upd)
);

/*Router 5,16*/    
cast_router #(
    .isUBM_list            (isUBM_list_5_16),
    .isFC_list             (isFC_list_5_16),
    .FCdn_list             (FCdn_list_5_16),
    .FCpl_list             (FCpl_list_5_16),
    .rt_file_list          (cast_rt_file_list_5_16)
)router_5_16(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_164_to_165),
    .west_valid_i          (valid_164_to_165),
    .west_ready_o          (ready_165_to_164),
    .west_data_o           (data_165_to_164),
    .west_valid_o          (valid_165_to_164),
    .west_ready_i          (ready_164_to_165),
    .east_data_i           (data_166_to_165),
    .east_valid_i          (valid_166_to_165),
    .east_ready_o          (ready_165_to_166),
    .east_data_o           (data_165_to_166),
    .east_valid_o          (valid_165_to_166),
    .east_ready_i          (ready_166_to_165),
    .vert0_data_i          (data_155_to_165_v0),
    .vert0_valid_i         (valid_155_to_165_v0),
    .vert0_ready_o         (ready_165_to_155_v0),
    .vert0_data_o          (data_165_to_175_v0),
    .vert0_valid_o         (valid_165_to_175_v0),
    .vert0_ready_i         (ready_175_to_165_v0),
    .vert1_data_i          (data_155_to_165_v1),
    .vert1_valid_i         (valid_155_to_165_v1),
    .vert1_ready_o         (ready_165_to_155_v1),
    .vert1_data_o          (data_165_to_175_v1),
    .vert1_valid_o         (valid_165_to_175_v1),
    .vert1_ready_i         (ready_175_to_165_v1),
    .local_data_i          (data_i[5][16]),
    .local_valid_i         (valid_i[5][16]),
    .local_ready_o         (ready_o[5][16]),
    .local_data_o          (data_o[5][16]),
    .local_valid_o         (valid_o[5][16]),
    .local_ready_i         (ready_i[5][16]),
    .credit_upd            (credit_upd)
);

/*Router 5,17*/    
cast_router #(
    .isUBM_list            (isUBM_list_5_17),
    .isFC_list             (isFC_list_5_17),
    .FCdn_list             (FCdn_list_5_17),
    .FCpl_list             (FCpl_list_5_17),
    .rt_file_list          (cast_rt_file_list_5_17)
)router_5_17(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_174_to_175),
    .west_valid_i          (valid_174_to_175),
    .west_ready_o          (ready_175_to_174),
    .west_data_o           (data_175_to_174),
    .west_valid_o          (valid_175_to_174),
    .west_ready_i          (ready_174_to_175),
    .east_data_i           (data_176_to_175),
    .east_valid_i          (valid_176_to_175),
    .east_ready_o          (ready_175_to_176),
    .east_data_o           (data_175_to_176),
    .east_valid_o          (valid_175_to_176),
    .east_ready_i          (ready_176_to_175),
    .vert0_data_i          (data_165_to_175_v0),
    .vert0_valid_i         (valid_165_to_175_v0),
    .vert0_ready_o         (ready_175_to_165_v0),
    .vert0_data_o          (data_175_to_185_v0),
    .vert0_valid_o         (valid_175_to_185_v0),
    .vert0_ready_i         (ready_185_to_175_v0),
    .vert1_data_i          (data_165_to_175_v1),
    .vert1_valid_i         (valid_165_to_175_v1),
    .vert1_ready_o         (ready_175_to_165_v1),
    .vert1_data_o          (data_175_to_185_v1),
    .vert1_valid_o         (valid_175_to_185_v1),
    .vert1_ready_i         (ready_185_to_175_v1),
    .local_data_i          (data_i[5][17]),
    .local_valid_i         (valid_i[5][17]),
    .local_ready_o         (ready_o[5][17]),
    .local_data_o          (data_o[5][17]),
    .local_valid_o         (valid_o[5][17]),
    .local_ready_i         (ready_i[5][17]),
    .credit_upd            (credit_upd)
);

/*Router 5,18*/    
cast_router #(
    .isUBM_list            (isUBM_list_5_18),
    .isFC_list             (isFC_list_5_18),
    .FCdn_list             (FCdn_list_5_18),
    .FCpl_list             (FCpl_list_5_18),
    .rt_file_list          (cast_rt_file_list_5_18)
)router_5_18(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_184_to_185),
    .west_valid_i          (valid_184_to_185),
    .west_ready_o          (ready_185_to_184),
    .west_data_o           (data_185_to_184),
    .west_valid_o          (valid_185_to_184),
    .west_ready_i          (ready_184_to_185),
    .east_data_i           (data_186_to_185),
    .east_valid_i          (valid_186_to_185),
    .east_ready_o          (ready_185_to_186),
    .east_data_o           (data_185_to_186),
    .east_valid_o          (valid_185_to_186),
    .east_ready_i          (ready_186_to_185),
    .vert0_data_i          (data_175_to_185_v0),
    .vert0_valid_i         (valid_175_to_185_v0),
    .vert0_ready_o         (ready_185_to_175_v0),
    .vert0_data_o          (data_185_to_195_v0),
    .vert0_valid_o         (valid_185_to_195_v0),
    .vert0_ready_i         (ready_195_to_185_v0),
    .vert1_data_i          (data_175_to_185_v1),
    .vert1_valid_i         (valid_175_to_185_v1),
    .vert1_ready_o         (ready_185_to_175_v1),
    .vert1_data_o          (data_185_to_195_v1),
    .vert1_valid_o         (valid_185_to_195_v1),
    .vert1_ready_i         (ready_195_to_185_v1),
    .local_data_i          (data_i[5][18]),
    .local_valid_i         (valid_i[5][18]),
    .local_ready_o         (ready_o[5][18]),
    .local_data_o          (data_o[5][18]),
    .local_valid_o         (valid_o[5][18]),
    .local_ready_i         (ready_i[5][18]),
    .credit_upd            (credit_upd)
);

/*Router 5,19*/    
cast_router #(
    .isUBM_list            (isUBM_list_5_19),
    .isFC_list             (isFC_list_5_19),
    .FCdn_list             (FCdn_list_5_19),
    .FCpl_list             (FCpl_list_5_19),
    .rt_file_list          (cast_rt_file_list_5_19)
)router_5_19(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_194_to_195),
    .west_valid_i          (valid_194_to_195),
    .west_ready_o          (ready_195_to_194),
    .west_data_o           (data_195_to_194),
    .west_valid_o          (valid_195_to_194),
    .west_ready_i          (ready_194_to_195),
    .east_data_i           (data_196_to_195),
    .east_valid_i          (valid_196_to_195),
    .east_ready_o          (ready_195_to_196),
    .east_data_o           (data_195_to_196),
    .east_valid_o          (valid_195_to_196),
    .east_ready_i          (ready_196_to_195),
    .vert0_data_i          (data_185_to_195_v0),
    .vert0_valid_i         (valid_185_to_195_v0),
    .vert0_ready_o         (ready_195_to_185_v0),
    .vert0_data_o          (data_195_to_205_v0),
    .vert0_valid_o         (valid_195_to_205_v0),
    .vert0_ready_i         (ready_205_to_195_v0),
    .vert1_data_i          (data_185_to_195_v1),
    .vert1_valid_i         (valid_185_to_195_v1),
    .vert1_ready_o         (ready_195_to_185_v1),
    .vert1_data_o          (data_195_to_205_v1),
    .vert1_valid_o         (valid_195_to_205_v1),
    .vert1_ready_i         (ready_205_to_195_v1),
    .local_data_i          (data_i[5][19]),
    .local_valid_i         (valid_i[5][19]),
    .local_ready_o         (ready_o[5][19]),
    .local_data_o          (data_o[5][19]),
    .local_valid_o         (valid_o[5][19]),
    .local_ready_i         (ready_i[5][19]),
    .credit_upd            (credit_upd)
);

/*Router 5,20*/    
cast_router #(
    .isUBM_list            (isUBM_list_5_20),
    .isFC_list             (isFC_list_5_20),
    .FCdn_list             (FCdn_list_5_20),
    .FCpl_list             (FCpl_list_5_20),
    .rt_file_list          (cast_rt_file_list_5_20)
)router_5_20(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_204_to_205),
    .west_valid_i          (valid_204_to_205),
    .west_ready_o          (ready_205_to_204),
    .west_data_o           (data_205_to_204),
    .west_valid_o          (valid_205_to_204),
    .west_ready_i          (ready_204_to_205),
    .east_data_i           (data_206_to_205),
    .east_valid_i          (valid_206_to_205),
    .east_ready_o          (ready_205_to_206),
    .east_data_o           (data_205_to_206),
    .east_valid_o          (valid_205_to_206),
    .east_ready_i          (ready_206_to_205),
    .vert0_data_i          (data_195_to_205_v0),
    .vert0_valid_i         (valid_195_to_205_v0),
    .vert0_ready_o         (ready_205_to_195_v0),
    .vert0_data_o          (data_205_to_215_v0),
    .vert0_valid_o         (valid_205_to_215_v0),
    .vert0_ready_i         (ready_215_to_205_v0),
    .vert1_data_i          (data_195_to_205_v1),
    .vert1_valid_i         (valid_195_to_205_v1),
    .vert1_ready_o         (ready_205_to_195_v1),
    .vert1_data_o          (data_205_to_215_v1),
    .vert1_valid_o         (valid_205_to_215_v1),
    .vert1_ready_i         (ready_215_to_205_v1),
    .local_data_i          (data_i[5][20]),
    .local_valid_i         (valid_i[5][20]),
    .local_ready_o         (ready_o[5][20]),
    .local_data_o          (data_o[5][20]),
    .local_valid_o         (valid_o[5][20]),
    .local_ready_i         (ready_i[5][20]),
    .credit_upd            (credit_upd)
);

/*Router 5,21*/    
cast_router #(
    .isUBM_list            (isUBM_list_5_21),
    .isFC_list             (isFC_list_5_21),
    .FCdn_list             (FCdn_list_5_21),
    .FCpl_list             (FCpl_list_5_21),
    .rt_file_list          (cast_rt_file_list_5_21)
)router_5_21(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_214_to_215),
    .west_valid_i          (valid_214_to_215),
    .west_ready_o          (ready_215_to_214),
    .west_data_o           (data_215_to_214),
    .west_valid_o          (valid_215_to_214),
    .west_ready_i          (ready_214_to_215),
    .east_data_i           (data_216_to_215),
    .east_valid_i          (valid_216_to_215),
    .east_ready_o          (ready_215_to_216),
    .east_data_o           (data_215_to_216),
    .east_valid_o          (valid_215_to_216),
    .east_ready_i          (ready_216_to_215),
    .vert0_data_i          (data_205_to_215_v0),
    .vert0_valid_i         (valid_205_to_215_v0),
    .vert0_ready_o         (ready_215_to_205_v0),
    .vert0_data_o          (data_215_to_225_v0),
    .vert0_valid_o         (valid_215_to_225_v0),
    .vert0_ready_i         (ready_225_to_215_v0),
    .vert1_data_i          (data_205_to_215_v1),
    .vert1_valid_i         (valid_205_to_215_v1),
    .vert1_ready_o         (ready_215_to_205_v1),
    .vert1_data_o          (data_215_to_225_v1),
    .vert1_valid_o         (valid_215_to_225_v1),
    .vert1_ready_i         (ready_225_to_215_v1),
    .local_data_i          (data_i[5][21]),
    .local_valid_i         (valid_i[5][21]),
    .local_ready_o         (ready_o[5][21]),
    .local_data_o          (data_o[5][21]),
    .local_valid_o         (valid_o[5][21]),
    .local_ready_i         (ready_i[5][21]),
    .credit_upd            (credit_upd)
);

/*Router 5,22*/    
cast_router #(
    .isUBM_list            (isUBM_list_5_22),
    .isFC_list             (isFC_list_5_22),
    .FCdn_list             (FCdn_list_5_22),
    .FCpl_list             (FCpl_list_5_22),
    .rt_file_list          (cast_rt_file_list_5_22)
)router_5_22(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_224_to_225),
    .west_valid_i          (valid_224_to_225),
    .west_ready_o          (ready_225_to_224),
    .west_data_o           (data_225_to_224),
    .west_valid_o          (valid_225_to_224),
    .west_ready_i          (ready_224_to_225),
    .east_data_i           (data_226_to_225),
    .east_valid_i          (valid_226_to_225),
    .east_ready_o          (ready_225_to_226),
    .east_data_o           (data_225_to_226),
    .east_valid_o          (valid_225_to_226),
    .east_ready_i          (ready_226_to_225),
    .vert0_data_i          (data_215_to_225_v0),
    .vert0_valid_i         (valid_215_to_225_v0),
    .vert0_ready_o         (ready_225_to_215_v0),
    .vert0_data_o          (data_225_to_235_v0),
    .vert0_valid_o         (valid_225_to_235_v0),
    .vert0_ready_i         (ready_235_to_225_v0),
    .vert1_data_i          (data_215_to_225_v1),
    .vert1_valid_i         (valid_215_to_225_v1),
    .vert1_ready_o         (ready_225_to_215_v1),
    .vert1_data_o          (data_225_to_235_v1),
    .vert1_valid_o         (valid_225_to_235_v1),
    .vert1_ready_i         (ready_235_to_225_v1),
    .local_data_i          (data_i[5][22]),
    .local_valid_i         (valid_i[5][22]),
    .local_ready_o         (ready_o[5][22]),
    .local_data_o          (data_o[5][22]),
    .local_valid_o         (valid_o[5][22]),
    .local_ready_i         (ready_i[5][22]),
    .credit_upd            (credit_upd)
);

/*Router 5,23*/    
cast_router #(
    .isUBM_list            (isUBM_list_5_23),
    .isFC_list             (isFC_list_5_23),
    .FCdn_list             (FCdn_list_5_23),
    .FCpl_list             (FCpl_list_5_23),
    .rt_file_list          (cast_rt_file_list_5_23)
)router_5_23(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_234_to_235),
    .west_valid_i          (valid_234_to_235),
    .west_ready_o          (ready_235_to_234),
    .west_data_o           (data_o_flee4),
    .west_valid_o          (valid_o_flee4),
    .west_ready_i          (ready_i_flee4),
    .east_data_i           (data_236_to_235),
    .east_valid_i          (valid_236_to_235),
    .east_ready_o          (ready_235_to_236),
    .east_data_o           (data_235_to_236),
    .east_valid_o          (valid_235_to_236),
    .east_ready_i          (ready_236_to_235),
    .vert0_data_i          (data_225_to_235_v0),
    .vert0_valid_i         (valid_225_to_235_v0),
    .vert0_ready_o         (ready_235_to_225_v0),
    .vert0_data_o          (data_235_to_245_v0),
    .vert0_valid_o         (valid_235_to_245_v0),
    .vert0_ready_i         (ready_245_to_235_v0),
    .vert1_data_i          (data_225_to_235_v1),
    .vert1_valid_i         (valid_225_to_235_v1),
    .vert1_ready_o         (ready_235_to_225_v1),
    .vert1_data_o          (data_235_to_245_v1),
    .vert1_valid_o         (valid_235_to_245_v1),
    .vert1_ready_i         (ready_245_to_235_v1),
    .local_data_i          (data_i[5][23]),
    .local_valid_i         (valid_i[5][23]),
    .local_ready_o         (ready_o[5][23]),
    .local_data_o          (data_o[5][23]),
    .local_valid_o         (valid_o[5][23]),
    .local_ready_i         (ready_i[5][23]),
    .credit_upd            (credit_upd)
);

/*Router 5,24*/    
cast_router #(
    .isUBM_list            (isUBM_list_5_24),
    .isFC_list             (isFC_list_5_24),
    .FCdn_list             (FCdn_list_5_24),
    .FCpl_list             (FCpl_list_5_24),
    .rt_file_list          (cast_rt_file_list_5_24)
)router_5_24(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_244_to_245),
    .west_valid_i          (valid_244_to_245),
    .west_ready_o          (ready_245_to_244),
    .west_data_o           (data_245_to_244),
    .west_valid_o          (valid_245_to_244),
    .west_ready_i          (ready_244_to_245),
    .east_data_i           (data_246_to_245),
    .east_valid_i          (valid_246_to_245),
    .east_ready_o          (ready_245_to_246),
    .east_data_o           (data_245_to_246),
    .east_valid_o          (valid_245_to_246),
    .east_ready_i          (ready_246_to_245),
    .vert0_data_i          (data_235_to_245_v0),
    .vert0_valid_i         (valid_235_to_245_v0),
    .vert0_ready_o         (ready_245_to_235_v0),
    .vert0_data_o          (),
    .vert0_valid_o         (),
    .vert0_ready_i         (1'b0),
    .vert1_data_i          (data_235_to_245_v1),
    .vert1_valid_i         (valid_235_to_245_v1),
    .vert1_ready_o         (ready_245_to_235_v1),
    .vert1_data_o          (),
    .vert1_valid_o         (),
    .vert1_ready_i         (1'b0),
    .local_data_i          (data_i[5][24]),
    .local_valid_i         (valid_i[5][24]),
    .local_ready_o         (ready_o[5][24]),
    .local_data_o          (data_o[5][24]),
    .local_valid_o         (valid_o[5][24]),
    .local_ready_i         (ready_i[5][24]),
    .credit_upd            (credit_upd)
);

/*Router 6,0*/    
cast_router #(
    .isUBM_list            (isUBM_list_6_0),
    .isFC_list             (isFC_list_6_0),
    .FCdn_list             (FCdn_list_6_0),
    .FCpl_list             (FCpl_list_6_0),
    .rt_file_list          (cast_rt_file_list_6_0)
)router_6_0(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_5_to_6),
    .west_valid_i          (valid_5_to_6),
    .west_ready_o          (ready_6_to_5),
    .west_data_o           (data_6_to_5),
    .west_valid_o          (valid_6_to_5),
    .west_ready_i          (ready_5_to_6),
    .east_data_i           (data_7_to_6),
    .east_valid_i          (valid_7_to_6),
    .east_ready_o          (ready_6_to_7),
    .east_data_o           (data_6_to_7),
    .east_valid_o          (valid_6_to_7),
    .east_ready_i          (ready_7_to_6),
    .vert0_data_i          (34'b0),
    .vert0_valid_i         (1'b0),
    .vert0_ready_o         (),
    .vert0_data_o          (data_6_to_16_v0),
    .vert0_valid_o         (valid_6_to_16_v0),
    .vert0_ready_i         (ready_16_to_6_v0),
    .vert1_data_i          (34'b0),
    .vert1_valid_i         (1'b0),
    .vert1_ready_o         (),
    .vert1_data_o          (data_6_to_16_v1),
    .vert1_valid_o         (valid_6_to_16_v1),
    .vert1_ready_i         (ready_16_to_6_v1),
    .local_data_i          (data_i[6][0]),
    .local_valid_i         (valid_i[6][0]),
    .local_ready_o         (ready_o[6][0]),
    .local_data_o          (data_o[6][0]),
    .local_valid_o         (valid_o[6][0]),
    .local_ready_i         (ready_i[6][0]),
    .credit_upd            (credit_upd)
);

/*Router 6,1*/    
cast_router #(
    .isUBM_list            (isUBM_list_6_1),
    .isFC_list             (isFC_list_6_1),
    .FCdn_list             (FCdn_list_6_1),
    .FCpl_list             (FCpl_list_6_1),
    .rt_file_list          (cast_rt_file_list_6_1)
)router_6_1(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_15_to_16),
    .west_valid_i          (valid_15_to_16),
    .west_ready_o          (ready_16_to_15),
    .west_data_o           (data_16_to_15),
    .west_valid_o          (valid_16_to_15),
    .west_ready_i          (ready_15_to_16),
    .east_data_i           (data_17_to_16),
    .east_valid_i          (valid_17_to_16),
    .east_ready_o          (ready_16_to_17),
    .east_data_o           (data_16_to_17),
    .east_valid_o          (valid_16_to_17),
    .east_ready_i          (ready_17_to_16),
    .vert0_data_i          (data_6_to_16_v0),
    .vert0_valid_i         (valid_6_to_16_v0),
    .vert0_ready_o         (ready_16_to_6_v0),
    .vert0_data_o          (data_16_to_26_v0),
    .vert0_valid_o         (valid_16_to_26_v0),
    .vert0_ready_i         (ready_26_to_16_v0),
    .vert1_data_i          (data_6_to_16_v1),
    .vert1_valid_i         (valid_6_to_16_v1),
    .vert1_ready_o         (ready_16_to_6_v1),
    .vert1_data_o          (data_16_to_26_v1),
    .vert1_valid_o         (valid_16_to_26_v1),
    .vert1_ready_i         (ready_26_to_16_v1),
    .local_data_i          (data_i[6][1]),
    .local_valid_i         (valid_i[6][1]),
    .local_ready_o         (ready_o[6][1]),
    .local_data_o          (data_o[6][1]),
    .local_valid_o         (valid_o[6][1]),
    .local_ready_i         (ready_i[6][1]),
    .credit_upd            (credit_upd)
);

/*Router 6,2*/    
cast_router #(
    .isUBM_list            (isUBM_list_6_2),
    .isFC_list             (isFC_list_6_2),
    .FCdn_list             (FCdn_list_6_2),
    .FCpl_list             (FCpl_list_6_2),
    .rt_file_list          (cast_rt_file_list_6_2)
)router_6_2(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_25_to_26),
    .west_valid_i          (valid_25_to_26),
    .west_ready_o          (ready_26_to_25),
    .west_data_o           (data_26_to_25),
    .west_valid_o          (valid_26_to_25),
    .west_ready_i          (ready_25_to_26),
    .east_data_i           (data_27_to_26),
    .east_valid_i          (valid_27_to_26),
    .east_ready_o          (ready_26_to_27),
    .east_data_o           (data_26_to_27),
    .east_valid_o          (valid_26_to_27),
    .east_ready_i          (ready_27_to_26),
    .vert0_data_i          (data_16_to_26_v0),
    .vert0_valid_i         (valid_16_to_26_v0),
    .vert0_ready_o         (ready_26_to_16_v0),
    .vert0_data_o          (data_26_to_36_v0),
    .vert0_valid_o         (valid_26_to_36_v0),
    .vert0_ready_i         (ready_36_to_26_v0),
    .vert1_data_i          (data_16_to_26_v1),
    .vert1_valid_i         (valid_16_to_26_v1),
    .vert1_ready_o         (ready_26_to_16_v1),
    .vert1_data_o          (data_26_to_36_v1),
    .vert1_valid_o         (valid_26_to_36_v1),
    .vert1_ready_i         (ready_36_to_26_v1),
    .local_data_i          (data_i[6][2]),
    .local_valid_i         (valid_i[6][2]),
    .local_ready_o         (ready_o[6][2]),
    .local_data_o          (data_o[6][2]),
    .local_valid_o         (valid_o[6][2]),
    .local_ready_i         (ready_i[6][2]),
    .credit_upd            (credit_upd)
);

/*Router 6,3*/    
cast_router #(
    .isUBM_list            (isUBM_list_6_3),
    .isFC_list             (isFC_list_6_3),
    .FCdn_list             (FCdn_list_6_3),
    .FCpl_list             (FCpl_list_6_3),
    .rt_file_list          (cast_rt_file_list_6_3)
)router_6_3(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_35_to_36),
    .west_valid_i          (valid_35_to_36),
    .west_ready_o          (ready_36_to_35),
    .west_data_o           (data_36_to_35),
    .west_valid_o          (valid_36_to_35),
    .west_ready_i          (ready_35_to_36),
    .east_data_i           (data_37_to_36),
    .east_valid_i          (valid_37_to_36),
    .east_ready_o          (ready_36_to_37),
    .east_data_o           (data_36_to_37),
    .east_valid_o          (valid_36_to_37),
    .east_ready_i          (ready_37_to_36),
    .vert0_data_i          (data_26_to_36_v0),
    .vert0_valid_i         (valid_26_to_36_v0),
    .vert0_ready_o         (ready_36_to_26_v0),
    .vert0_data_o          (data_36_to_46_v0),
    .vert0_valid_o         (valid_36_to_46_v0),
    .vert0_ready_i         (ready_46_to_36_v0),
    .vert1_data_i          (data_26_to_36_v1),
    .vert1_valid_i         (valid_26_to_36_v1),
    .vert1_ready_o         (ready_36_to_26_v1),
    .vert1_data_o          (data_36_to_46_v1),
    .vert1_valid_o         (valid_36_to_46_v1),
    .vert1_ready_i         (ready_46_to_36_v1),
    .local_data_i          (data_i[6][3]),
    .local_valid_i         (valid_i[6][3]),
    .local_ready_o         (ready_o[6][3]),
    .local_data_o          (data_o[6][3]),
    .local_valid_o         (valid_o[6][3]),
    .local_ready_i         (ready_i[6][3]),
    .credit_upd            (credit_upd)
);

/*Router 6,4*/    
cast_router #(
    .isUBM_list            (isUBM_list_6_4),
    .isFC_list             (isFC_list_6_4),
    .FCdn_list             (FCdn_list_6_4),
    .FCpl_list             (FCpl_list_6_4),
    .rt_file_list          (cast_rt_file_list_6_4)
)router_6_4(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_45_to_46),
    .west_valid_i          (valid_45_to_46),
    .west_ready_o          (ready_46_to_45),
    .west_data_o           (data_46_to_45),
    .west_valid_o          (valid_46_to_45),
    .west_ready_i          (ready_45_to_46),
    .east_data_i           (data_47_to_46),
    .east_valid_i          (valid_47_to_46),
    .east_ready_o          (ready_46_to_47),
    .east_data_o           (data_46_to_47),
    .east_valid_o          (valid_46_to_47),
    .east_ready_i          (ready_47_to_46),
    .vert0_data_i          (data_36_to_46_v0),
    .vert0_valid_i         (valid_36_to_46_v0),
    .vert0_ready_o         (ready_46_to_36_v0),
    .vert0_data_o          (data_46_to_56_v0),
    .vert0_valid_o         (valid_46_to_56_v0),
    .vert0_ready_i         (ready_56_to_46_v0),
    .vert1_data_i          (data_36_to_46_v1),
    .vert1_valid_i         (valid_36_to_46_v1),
    .vert1_ready_o         (ready_46_to_36_v1),
    .vert1_data_o          (data_46_to_56_v1),
    .vert1_valid_o         (valid_46_to_56_v1),
    .vert1_ready_i         (ready_56_to_46_v1),
    .local_data_i          (data_i[6][4]),
    .local_valid_i         (valid_i[6][4]),
    .local_ready_o         (ready_o[6][4]),
    .local_data_o          (data_o[6][4]),
    .local_valid_o         (valid_o[6][4]),
    .local_ready_i         (ready_i[6][4]),
    .credit_upd            (credit_upd)
);

/*Router 6,5*/    
cast_router #(
    .isUBM_list            (isUBM_list_6_5),
    .isFC_list             (isFC_list_6_5),
    .FCdn_list             (FCdn_list_6_5),
    .FCpl_list             (FCpl_list_6_5),
    .rt_file_list          (cast_rt_file_list_6_5)
)router_6_5(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_55_to_56),
    .west_valid_i          (valid_55_to_56),
    .west_ready_o          (ready_56_to_55),
    .west_data_o           (data_56_to_55),
    .west_valid_o          (valid_56_to_55),
    .west_ready_i          (ready_55_to_56),
    .east_data_i           (data_57_to_56),
    .east_valid_i          (valid_57_to_56),
    .east_ready_o          (ready_56_to_57),
    .east_data_o           (data_56_to_57),
    .east_valid_o          (valid_56_to_57),
    .east_ready_i          (ready_57_to_56),
    .vert0_data_i          (data_46_to_56_v0),
    .vert0_valid_i         (valid_46_to_56_v0),
    .vert0_ready_o         (ready_56_to_46_v0),
    .vert0_data_o          (data_56_to_66_v0),
    .vert0_valid_o         (valid_56_to_66_v0),
    .vert0_ready_i         (ready_66_to_56_v0),
    .vert1_data_i          (data_46_to_56_v1),
    .vert1_valid_i         (valid_46_to_56_v1),
    .vert1_ready_o         (ready_56_to_46_v1),
    .vert1_data_o          (data_56_to_66_v1),
    .vert1_valid_o         (valid_56_to_66_v1),
    .vert1_ready_i         (ready_66_to_56_v1),
    .local_data_i          (data_i[6][5]),
    .local_valid_i         (valid_i[6][5]),
    .local_ready_o         (ready_o[6][5]),
    .local_data_o          (data_o[6][5]),
    .local_valid_o         (valid_o[6][5]),
    .local_ready_i         (ready_i[6][5]),
    .credit_upd            (credit_upd)
);

/*Router 6,6*/    
cast_router #(
    .isUBM_list            (isUBM_list_6_6),
    .isFC_list             (isFC_list_6_6),
    .FCdn_list             (FCdn_list_6_6),
    .FCpl_list             (FCpl_list_6_6),
    .rt_file_list          (cast_rt_file_list_6_6)
)router_6_6(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_65_to_66),
    .west_valid_i          (valid_65_to_66),
    .west_ready_o          (ready_66_to_65),
    .west_data_o           (data_66_to_65),
    .west_valid_o          (valid_66_to_65),
    .west_ready_i          (ready_65_to_66),
    .east_data_i           (data_67_to_66),
    .east_valid_i          (valid_67_to_66),
    .east_ready_o          (ready_66_to_67),
    .east_data_o           (data_66_to_67),
    .east_valid_o          (valid_66_to_67),
    .east_ready_i          (ready_67_to_66),
    .vert0_data_i          (data_56_to_66_v0),
    .vert0_valid_i         (valid_56_to_66_v0),
    .vert0_ready_o         (ready_66_to_56_v0),
    .vert0_data_o          (data_66_to_76_v0),
    .vert0_valid_o         (valid_66_to_76_v0),
    .vert0_ready_i         (ready_76_to_66_v0),
    .vert1_data_i          (data_56_to_66_v1),
    .vert1_valid_i         (valid_56_to_66_v1),
    .vert1_ready_o         (ready_66_to_56_v1),
    .vert1_data_o          (data_66_to_76_v1),
    .vert1_valid_o         (valid_66_to_76_v1),
    .vert1_ready_i         (ready_76_to_66_v1),
    .local_data_i          (data_i[6][6]),
    .local_valid_i         (valid_i[6][6]),
    .local_ready_o         (ready_o[6][6]),
    .local_data_o          (data_o[6][6]),
    .local_valid_o         (valid_o[6][6]),
    .local_ready_i         (ready_i[6][6]),
    .credit_upd            (credit_upd)
);

/*Router 6,7*/    
cast_router #(
    .isUBM_list            (isUBM_list_6_7),
    .isFC_list             (isFC_list_6_7),
    .FCdn_list             (FCdn_list_6_7),
    .FCpl_list             (FCpl_list_6_7),
    .rt_file_list          (cast_rt_file_list_6_7)
)router_6_7(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_75_to_76),
    .west_valid_i          (valid_75_to_76),
    .west_ready_o          (ready_76_to_75),
    .west_data_o           (data_76_to_75),
    .west_valid_o          (valid_76_to_75),
    .west_ready_i          (ready_75_to_76),
    .east_data_i           (data_77_to_76),
    .east_valid_i          (valid_77_to_76),
    .east_ready_o          (ready_76_to_77),
    .east_data_o           (data_76_to_77),
    .east_valid_o          (valid_76_to_77),
    .east_ready_i          (ready_77_to_76),
    .vert0_data_i          (data_66_to_76_v0),
    .vert0_valid_i         (valid_66_to_76_v0),
    .vert0_ready_o         (ready_76_to_66_v0),
    .vert0_data_o          (data_76_to_86_v0),
    .vert0_valid_o         (valid_76_to_86_v0),
    .vert0_ready_i         (ready_86_to_76_v0),
    .vert1_data_i          (data_66_to_76_v1),
    .vert1_valid_i         (valid_66_to_76_v1),
    .vert1_ready_o         (ready_76_to_66_v1),
    .vert1_data_o          (data_76_to_86_v1),
    .vert1_valid_o         (valid_76_to_86_v1),
    .vert1_ready_i         (ready_86_to_76_v1),
    .local_data_i          (data_i[6][7]),
    .local_valid_i         (valid_i[6][7]),
    .local_ready_o         (ready_o[6][7]),
    .local_data_o          (data_o[6][7]),
    .local_valid_o         (valid_o[6][7]),
    .local_ready_i         (ready_i[6][7]),
    .credit_upd            (credit_upd)
);

/*Router 6,8*/    
cast_router #(
    .isUBM_list            (isUBM_list_6_8),
    .isFC_list             (isFC_list_6_8),
    .FCdn_list             (FCdn_list_6_8),
    .FCpl_list             (FCpl_list_6_8),
    .rt_file_list          (cast_rt_file_list_6_8)
)router_6_8(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_85_to_86),
    .west_valid_i          (valid_85_to_86),
    .west_ready_o          (ready_86_to_85),
    .west_data_o           (data_86_to_85),
    .west_valid_o          (valid_86_to_85),
    .west_ready_i          (ready_85_to_86),
    .east_data_i           (data_87_to_86),
    .east_valid_i          (valid_87_to_86),
    .east_ready_o          (ready_86_to_87),
    .east_data_o           (data_86_to_87),
    .east_valid_o          (valid_86_to_87),
    .east_ready_i          (ready_87_to_86),
    .vert0_data_i          (data_76_to_86_v0),
    .vert0_valid_i         (valid_76_to_86_v0),
    .vert0_ready_o         (ready_86_to_76_v0),
    .vert0_data_o          (data_86_to_96_v0),
    .vert0_valid_o         (valid_86_to_96_v0),
    .vert0_ready_i         (ready_96_to_86_v0),
    .vert1_data_i          (data_76_to_86_v1),
    .vert1_valid_i         (valid_76_to_86_v1),
    .vert1_ready_o         (ready_86_to_76_v1),
    .vert1_data_o          (data_86_to_96_v1),
    .vert1_valid_o         (valid_86_to_96_v1),
    .vert1_ready_i         (ready_96_to_86_v1),
    .local_data_i          (data_i[6][8]),
    .local_valid_i         (valid_i[6][8]),
    .local_ready_o         (ready_o[6][8]),
    .local_data_o          (data_o[6][8]),
    .local_valid_o         (valid_o[6][8]),
    .local_ready_i         (ready_i[6][8]),
    .credit_upd            (credit_upd)
);

/*Router 6,9*/    
cast_router #(
    .isUBM_list            (isUBM_list_6_9),
    .isFC_list             (isFC_list_6_9),
    .FCdn_list             (FCdn_list_6_9),
    .FCpl_list             (FCpl_list_6_9),
    .rt_file_list          (cast_rt_file_list_6_9)
)router_6_9(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_95_to_96),
    .west_valid_i          (valid_95_to_96),
    .west_ready_o          (ready_96_to_95),
    .west_data_o           (data_96_to_95),
    .west_valid_o          (valid_96_to_95),
    .west_ready_i          (ready_95_to_96),
    .east_data_i           (data_97_to_96),
    .east_valid_i          (valid_97_to_96),
    .east_ready_o          (ready_96_to_97),
    .east_data_o           (data_96_to_97),
    .east_valid_o          (valid_96_to_97),
    .east_ready_i          (ready_97_to_96),
    .vert0_data_i          (data_86_to_96_v0),
    .vert0_valid_i         (valid_86_to_96_v0),
    .vert0_ready_o         (ready_96_to_86_v0),
    .vert0_data_o          (data_96_to_106_v0),
    .vert0_valid_o         (valid_96_to_106_v0),
    .vert0_ready_i         (ready_106_to_96_v0),
    .vert1_data_i          (data_86_to_96_v1),
    .vert1_valid_i         (valid_86_to_96_v1),
    .vert1_ready_o         (ready_96_to_86_v1),
    .vert1_data_o          (data_96_to_106_v1),
    .vert1_valid_o         (valid_96_to_106_v1),
    .vert1_ready_i         (ready_106_to_96_v1),
    .local_data_i          (data_i[6][9]),
    .local_valid_i         (valid_i[6][9]),
    .local_ready_o         (ready_o[6][9]),
    .local_data_o          (data_o[6][9]),
    .local_valid_o         (valid_o[6][9]),
    .local_ready_i         (ready_i[6][9]),
    .credit_upd            (credit_upd)
);

/*Router 6,10*/    
cast_router #(
    .isUBM_list            (isUBM_list_6_10),
    .isFC_list             (isFC_list_6_10),
    .FCdn_list             (FCdn_list_6_10),
    .FCpl_list             (FCpl_list_6_10),
    .rt_file_list          (cast_rt_file_list_6_10)
)router_6_10(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_105_to_106),
    .west_valid_i          (valid_105_to_106),
    .west_ready_o          (ready_106_to_105),
    .west_data_o           (data_106_to_105),
    .west_valid_o          (valid_106_to_105),
    .west_ready_i          (ready_105_to_106),
    .east_data_i           (data_107_to_106),
    .east_valid_i          (valid_107_to_106),
    .east_ready_o          (ready_106_to_107),
    .east_data_o           (data_106_to_107),
    .east_valid_o          (valid_106_to_107),
    .east_ready_i          (ready_107_to_106),
    .vert0_data_i          (data_96_to_106_v0),
    .vert0_valid_i         (valid_96_to_106_v0),
    .vert0_ready_o         (ready_106_to_96_v0),
    .vert0_data_o          (data_106_to_116_v0),
    .vert0_valid_o         (valid_106_to_116_v0),
    .vert0_ready_i         (ready_116_to_106_v0),
    .vert1_data_i          (data_96_to_106_v1),
    .vert1_valid_i         (valid_96_to_106_v1),
    .vert1_ready_o         (ready_106_to_96_v1),
    .vert1_data_o          (data_106_to_116_v1),
    .vert1_valid_o         (valid_106_to_116_v1),
    .vert1_ready_i         (ready_116_to_106_v1),
    .local_data_i          (data_i[6][10]),
    .local_valid_i         (valid_i[6][10]),
    .local_ready_o         (ready_o[6][10]),
    .local_data_o          (data_o[6][10]),
    .local_valid_o         (valid_o[6][10]),
    .local_ready_i         (ready_i[6][10]),
    .credit_upd            (credit_upd)
);

/*Router 6,11*/    
cast_router #(
    .isUBM_list            (isUBM_list_6_11),
    .isFC_list             (isFC_list_6_11),
    .FCdn_list             (FCdn_list_6_11),
    .FCpl_list             (FCpl_list_6_11),
    .rt_file_list          (cast_rt_file_list_6_11)
)router_6_11(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_115_to_116),
    .west_valid_i          (valid_115_to_116),
    .west_ready_o          (ready_116_to_115),
    .west_data_o           (data_116_to_115),
    .west_valid_o          (valid_116_to_115),
    .west_ready_i          (ready_115_to_116),
    .east_data_i           (data_117_to_116),
    .east_valid_i          (valid_117_to_116),
    .east_ready_o          (ready_116_to_117),
    .east_data_o           (data_116_to_117),
    .east_valid_o          (valid_116_to_117),
    .east_ready_i          (ready_117_to_116),
    .vert0_data_i          (data_106_to_116_v0),
    .vert0_valid_i         (valid_106_to_116_v0),
    .vert0_ready_o         (ready_116_to_106_v0),
    .vert0_data_o          (data_116_to_126_v0),
    .vert0_valid_o         (valid_116_to_126_v0),
    .vert0_ready_i         (ready_126_to_116_v0),
    .vert1_data_i          (data_106_to_116_v1),
    .vert1_valid_i         (valid_106_to_116_v1),
    .vert1_ready_o         (ready_116_to_106_v1),
    .vert1_data_o          (data_116_to_126_v1),
    .vert1_valid_o         (valid_116_to_126_v1),
    .vert1_ready_i         (ready_126_to_116_v1),
    .local_data_i          (data_i[6][11]),
    .local_valid_i         (valid_i[6][11]),
    .local_ready_o         (ready_o[6][11]),
    .local_data_o          (data_o[6][11]),
    .local_valid_o         (valid_o[6][11]),
    .local_ready_i         (ready_i[6][11]),
    .credit_upd            (credit_upd)
);

/*Router 6,12*/    
cast_router #(
    .isUBM_list            (isUBM_list_6_12),
    .isFC_list             (isFC_list_6_12),
    .FCdn_list             (FCdn_list_6_12),
    .FCpl_list             (FCpl_list_6_12),
    .rt_file_list          (cast_rt_file_list_6_12)
)router_6_12(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_125_to_126),
    .west_valid_i          (valid_125_to_126),
    .west_ready_o          (ready_126_to_125),
    .west_data_o           (data_126_to_125),
    .west_valid_o          (valid_126_to_125),
    .west_ready_i          (ready_125_to_126),
    .east_data_i           (data_127_to_126),
    .east_valid_i          (valid_127_to_126),
    .east_ready_o          (ready_126_to_127),
    .east_data_o           (data_126_to_127),
    .east_valid_o          (valid_126_to_127),
    .east_ready_i          (ready_127_to_126),
    .vert0_data_i          (data_116_to_126_v0),
    .vert0_valid_i         (valid_116_to_126_v0),
    .vert0_ready_o         (ready_126_to_116_v0),
    .vert0_data_o          (data_126_to_136_v0),
    .vert0_valid_o         (valid_126_to_136_v0),
    .vert0_ready_i         (ready_136_to_126_v0),
    .vert1_data_i          (data_116_to_126_v1),
    .vert1_valid_i         (valid_116_to_126_v1),
    .vert1_ready_o         (ready_126_to_116_v1),
    .vert1_data_o          (data_126_to_136_v1),
    .vert1_valid_o         (valid_126_to_136_v1),
    .vert1_ready_i         (ready_136_to_126_v1),
    .local_data_i          (data_i[6][12]),
    .local_valid_i         (valid_i[6][12]),
    .local_ready_o         (ready_o[6][12]),
    .local_data_o          (data_o[6][12]),
    .local_valid_o         (valid_o[6][12]),
    .local_ready_i         (ready_i[6][12]),
    .credit_upd            (credit_upd)
);

/*Router 6,13*/    
cast_router #(
    .isUBM_list            (isUBM_list_6_13),
    .isFC_list             (isFC_list_6_13),
    .FCdn_list             (FCdn_list_6_13),
    .FCpl_list             (FCpl_list_6_13),
    .rt_file_list          (cast_rt_file_list_6_13)
)router_6_13(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_135_to_136),
    .west_valid_i          (valid_135_to_136),
    .west_ready_o          (ready_136_to_135),
    .west_data_o           (data_136_to_135),
    .west_valid_o          (valid_136_to_135),
    .west_ready_i          (ready_135_to_136),
    .east_data_i           (data_137_to_136),
    .east_valid_i          (valid_137_to_136),
    .east_ready_o          (ready_136_to_137),
    .east_data_o           (data_136_to_137),
    .east_valid_o          (valid_136_to_137),
    .east_ready_i          (ready_137_to_136),
    .vert0_data_i          (data_126_to_136_v0),
    .vert0_valid_i         (valid_126_to_136_v0),
    .vert0_ready_o         (ready_136_to_126_v0),
    .vert0_data_o          (data_136_to_146_v0),
    .vert0_valid_o         (valid_136_to_146_v0),
    .vert0_ready_i         (ready_146_to_136_v0),
    .vert1_data_i          (data_126_to_136_v1),
    .vert1_valid_i         (valid_126_to_136_v1),
    .vert1_ready_o         (ready_136_to_126_v1),
    .vert1_data_o          (data_136_to_146_v1),
    .vert1_valid_o         (valid_136_to_146_v1),
    .vert1_ready_i         (ready_146_to_136_v1),
    .local_data_i          (data_i[6][13]),
    .local_valid_i         (valid_i[6][13]),
    .local_ready_o         (ready_o[6][13]),
    .local_data_o          (data_o[6][13]),
    .local_valid_o         (valid_o[6][13]),
    .local_ready_i         (ready_i[6][13]),
    .credit_upd            (credit_upd)
);

/*Router 6,14*/    
cast_router #(
    .isUBM_list            (isUBM_list_6_14),
    .isFC_list             (isFC_list_6_14),
    .FCdn_list             (FCdn_list_6_14),
    .FCpl_list             (FCpl_list_6_14),
    .rt_file_list          (cast_rt_file_list_6_14)
)router_6_14(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_145_to_146),
    .west_valid_i          (valid_145_to_146),
    .west_ready_o          (ready_146_to_145),
    .west_data_o           (data_146_to_145),
    .west_valid_o          (valid_146_to_145),
    .west_ready_i          (ready_145_to_146),
    .east_data_i           (data_147_to_146),
    .east_valid_i          (valid_147_to_146),
    .east_ready_o          (ready_146_to_147),
    .east_data_o           (data_146_to_147),
    .east_valid_o          (valid_146_to_147),
    .east_ready_i          (ready_147_to_146),
    .vert0_data_i          (data_136_to_146_v0),
    .vert0_valid_i         (valid_136_to_146_v0),
    .vert0_ready_o         (ready_146_to_136_v0),
    .vert0_data_o          (data_146_to_156_v0),
    .vert0_valid_o         (valid_146_to_156_v0),
    .vert0_ready_i         (ready_156_to_146_v0),
    .vert1_data_i          (data_136_to_146_v1),
    .vert1_valid_i         (valid_136_to_146_v1),
    .vert1_ready_o         (ready_146_to_136_v1),
    .vert1_data_o          (data_146_to_156_v1),
    .vert1_valid_o         (valid_146_to_156_v1),
    .vert1_ready_i         (ready_156_to_146_v1),
    .local_data_i          (data_i[6][14]),
    .local_valid_i         (valid_i[6][14]),
    .local_ready_o         (ready_o[6][14]),
    .local_data_o          (data_o[6][14]),
    .local_valid_o         (valid_o[6][14]),
    .local_ready_i         (ready_i[6][14]),
    .credit_upd            (credit_upd)
);

/*Router 6,15*/    
cast_router #(
    .isUBM_list            (isUBM_list_6_15),
    .isFC_list             (isFC_list_6_15),
    .FCdn_list             (FCdn_list_6_15),
    .FCpl_list             (FCpl_list_6_15),
    .rt_file_list          (cast_rt_file_list_6_15)
)router_6_15(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_155_to_156),
    .west_valid_i          (valid_155_to_156),
    .west_ready_o          (ready_156_to_155),
    .west_data_o           (data_156_to_155),
    .west_valid_o          (valid_156_to_155),
    .west_ready_i          (ready_155_to_156),
    .east_data_i           (data_157_to_156),
    .east_valid_i          (valid_157_to_156),
    .east_ready_o          (ready_156_to_157),
    .east_data_o           (data_156_to_157),
    .east_valid_o          (valid_156_to_157),
    .east_ready_i          (ready_157_to_156),
    .vert0_data_i          (data_146_to_156_v0),
    .vert0_valid_i         (valid_146_to_156_v0),
    .vert0_ready_o         (ready_156_to_146_v0),
    .vert0_data_o          (data_156_to_166_v0),
    .vert0_valid_o         (valid_156_to_166_v0),
    .vert0_ready_i         (ready_166_to_156_v0),
    .vert1_data_i          (data_146_to_156_v1),
    .vert1_valid_i         (valid_146_to_156_v1),
    .vert1_ready_o         (ready_156_to_146_v1),
    .vert1_data_o          (data_156_to_166_v1),
    .vert1_valid_o         (valid_156_to_166_v1),
    .vert1_ready_i         (ready_166_to_156_v1),
    .local_data_i          (data_i[6][15]),
    .local_valid_i         (valid_i[6][15]),
    .local_ready_o         (ready_o[6][15]),
    .local_data_o          (data_o[6][15]),
    .local_valid_o         (valid_o[6][15]),
    .local_ready_i         (ready_i[6][15]),
    .credit_upd            (credit_upd)
);

/*Router 6,16*/    
cast_router #(
    .isUBM_list            (isUBM_list_6_16),
    .isFC_list             (isFC_list_6_16),
    .FCdn_list             (FCdn_list_6_16),
    .FCpl_list             (FCpl_list_6_16),
    .rt_file_list          (cast_rt_file_list_6_16)
)router_6_16(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_165_to_166),
    .west_valid_i          (valid_165_to_166),
    .west_ready_o          (ready_166_to_165),
    .west_data_o           (data_166_to_165),
    .west_valid_o          (valid_166_to_165),
    .west_ready_i          (ready_165_to_166),
    .east_data_i           (data_167_to_166),
    .east_valid_i          (valid_167_to_166),
    .east_ready_o          (ready_166_to_167),
    .east_data_o           (data_166_to_167),
    .east_valid_o          (valid_166_to_167),
    .east_ready_i          (ready_167_to_166),
    .vert0_data_i          (data_156_to_166_v0),
    .vert0_valid_i         (valid_156_to_166_v0),
    .vert0_ready_o         (ready_166_to_156_v0),
    .vert0_data_o          (data_166_to_176_v0),
    .vert0_valid_o         (valid_166_to_176_v0),
    .vert0_ready_i         (ready_176_to_166_v0),
    .vert1_data_i          (data_156_to_166_v1),
    .vert1_valid_i         (valid_156_to_166_v1),
    .vert1_ready_o         (ready_166_to_156_v1),
    .vert1_data_o          (data_166_to_176_v1),
    .vert1_valid_o         (valid_166_to_176_v1),
    .vert1_ready_i         (ready_176_to_166_v1),
    .local_data_i          (data_i[6][16]),
    .local_valid_i         (valid_i[6][16]),
    .local_ready_o         (ready_o[6][16]),
    .local_data_o          (data_o[6][16]),
    .local_valid_o         (valid_o[6][16]),
    .local_ready_i         (ready_i[6][16]),
    .credit_upd            (credit_upd)
);

/*Router 6,17*/    
cast_router #(
    .isUBM_list            (isUBM_list_6_17),
    .isFC_list             (isFC_list_6_17),
    .FCdn_list             (FCdn_list_6_17),
    .FCpl_list             (FCpl_list_6_17),
    .rt_file_list          (cast_rt_file_list_6_17)
)router_6_17(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_175_to_176),
    .west_valid_i          (valid_175_to_176),
    .west_ready_o          (ready_176_to_175),
    .west_data_o           (data_176_to_175),
    .west_valid_o          (valid_176_to_175),
    .west_ready_i          (ready_175_to_176),
    .east_data_i           (data_177_to_176),
    .east_valid_i          (valid_177_to_176),
    .east_ready_o          (ready_176_to_177),
    .east_data_o           (data_176_to_177),
    .east_valid_o          (valid_176_to_177),
    .east_ready_i          (ready_177_to_176),
    .vert0_data_i          (data_166_to_176_v0),
    .vert0_valid_i         (valid_166_to_176_v0),
    .vert0_ready_o         (ready_176_to_166_v0),
    .vert0_data_o          (data_176_to_186_v0),
    .vert0_valid_o         (valid_176_to_186_v0),
    .vert0_ready_i         (ready_186_to_176_v0),
    .vert1_data_i          (data_166_to_176_v1),
    .vert1_valid_i         (valid_166_to_176_v1),
    .vert1_ready_o         (ready_176_to_166_v1),
    .vert1_data_o          (data_176_to_186_v1),
    .vert1_valid_o         (valid_176_to_186_v1),
    .vert1_ready_i         (ready_186_to_176_v1),
    .local_data_i          (data_i[6][17]),
    .local_valid_i         (valid_i[6][17]),
    .local_ready_o         (ready_o[6][17]),
    .local_data_o          (data_o[6][17]),
    .local_valid_o         (valid_o[6][17]),
    .local_ready_i         (ready_i[6][17]),
    .credit_upd            (credit_upd)
);

/*Router 6,18*/    
cast_router #(
    .isUBM_list            (isUBM_list_6_18),
    .isFC_list             (isFC_list_6_18),
    .FCdn_list             (FCdn_list_6_18),
    .FCpl_list             (FCpl_list_6_18),
    .rt_file_list          (cast_rt_file_list_6_18)
)router_6_18(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_185_to_186),
    .west_valid_i          (valid_185_to_186),
    .west_ready_o          (ready_186_to_185),
    .west_data_o           (data_186_to_185),
    .west_valid_o          (valid_186_to_185),
    .west_ready_i          (ready_185_to_186),
    .east_data_i           (data_187_to_186),
    .east_valid_i          (valid_187_to_186),
    .east_ready_o          (ready_186_to_187),
    .east_data_o           (data_186_to_187),
    .east_valid_o          (valid_186_to_187),
    .east_ready_i          (ready_187_to_186),
    .vert0_data_i          (data_176_to_186_v0),
    .vert0_valid_i         (valid_176_to_186_v0),
    .vert0_ready_o         (ready_186_to_176_v0),
    .vert0_data_o          (data_186_to_196_v0),
    .vert0_valid_o         (valid_186_to_196_v0),
    .vert0_ready_i         (ready_196_to_186_v0),
    .vert1_data_i          (data_176_to_186_v1),
    .vert1_valid_i         (valid_176_to_186_v1),
    .vert1_ready_o         (ready_186_to_176_v1),
    .vert1_data_o          (data_186_to_196_v1),
    .vert1_valid_o         (valid_186_to_196_v1),
    .vert1_ready_i         (ready_196_to_186_v1),
    .local_data_i          (data_i[6][18]),
    .local_valid_i         (valid_i[6][18]),
    .local_ready_o         (ready_o[6][18]),
    .local_data_o          (data_o[6][18]),
    .local_valid_o         (valid_o[6][18]),
    .local_ready_i         (ready_i[6][18]),
    .credit_upd            (credit_upd)
);

/*Router 6,19*/    
cast_router #(
    .isUBM_list            (isUBM_list_6_19),
    .isFC_list             (isFC_list_6_19),
    .FCdn_list             (FCdn_list_6_19),
    .FCpl_list             (FCpl_list_6_19),
    .rt_file_list          (cast_rt_file_list_6_19)
)router_6_19(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_195_to_196),
    .west_valid_i          (valid_195_to_196),
    .west_ready_o          (ready_196_to_195),
    .west_data_o           (data_196_to_195),
    .west_valid_o          (valid_196_to_195),
    .west_ready_i          (ready_195_to_196),
    .east_data_i           (data_197_to_196),
    .east_valid_i          (valid_197_to_196),
    .east_ready_o          (ready_196_to_197),
    .east_data_o           (data_196_to_197),
    .east_valid_o          (valid_196_to_197),
    .east_ready_i          (ready_197_to_196),
    .vert0_data_i          (data_186_to_196_v0),
    .vert0_valid_i         (valid_186_to_196_v0),
    .vert0_ready_o         (ready_196_to_186_v0),
    .vert0_data_o          (data_196_to_206_v0),
    .vert0_valid_o         (valid_196_to_206_v0),
    .vert0_ready_i         (ready_206_to_196_v0),
    .vert1_data_i          (data_186_to_196_v1),
    .vert1_valid_i         (valid_186_to_196_v1),
    .vert1_ready_o         (ready_196_to_186_v1),
    .vert1_data_o          (data_196_to_206_v1),
    .vert1_valid_o         (valid_196_to_206_v1),
    .vert1_ready_i         (ready_206_to_196_v1),
    .local_data_i          (data_i[6][19]),
    .local_valid_i         (valid_i[6][19]),
    .local_ready_o         (ready_o[6][19]),
    .local_data_o          (data_o[6][19]),
    .local_valid_o         (valid_o[6][19]),
    .local_ready_i         (ready_i[6][19]),
    .credit_upd            (credit_upd)
);

/*Router 6,20*/    
cast_router #(
    .isUBM_list            (isUBM_list_6_20),
    .isFC_list             (isFC_list_6_20),
    .FCdn_list             (FCdn_list_6_20),
    .FCpl_list             (FCpl_list_6_20),
    .rt_file_list          (cast_rt_file_list_6_20)
)router_6_20(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_205_to_206),
    .west_valid_i          (valid_205_to_206),
    .west_ready_o          (ready_206_to_205),
    .west_data_o           (data_206_to_205),
    .west_valid_o          (valid_206_to_205),
    .west_ready_i          (ready_205_to_206),
    .east_data_i           (data_207_to_206),
    .east_valid_i          (valid_207_to_206),
    .east_ready_o          (ready_206_to_207),
    .east_data_o           (data_206_to_207),
    .east_valid_o          (valid_206_to_207),
    .east_ready_i          (ready_207_to_206),
    .vert0_data_i          (data_196_to_206_v0),
    .vert0_valid_i         (valid_196_to_206_v0),
    .vert0_ready_o         (ready_206_to_196_v0),
    .vert0_data_o          (data_206_to_216_v0),
    .vert0_valid_o         (valid_206_to_216_v0),
    .vert0_ready_i         (ready_216_to_206_v0),
    .vert1_data_i          (data_196_to_206_v1),
    .vert1_valid_i         (valid_196_to_206_v1),
    .vert1_ready_o         (ready_206_to_196_v1),
    .vert1_data_o          (data_206_to_216_v1),
    .vert1_valid_o         (valid_206_to_216_v1),
    .vert1_ready_i         (ready_216_to_206_v1),
    .local_data_i          (data_i[6][20]),
    .local_valid_i         (valid_i[6][20]),
    .local_ready_o         (ready_o[6][20]),
    .local_data_o          (data_o[6][20]),
    .local_valid_o         (valid_o[6][20]),
    .local_ready_i         (ready_i[6][20]),
    .credit_upd            (credit_upd)
);

/*Router 6,21*/    
cast_router #(
    .isUBM_list            (isUBM_list_6_21),
    .isFC_list             (isFC_list_6_21),
    .FCdn_list             (FCdn_list_6_21),
    .FCpl_list             (FCpl_list_6_21),
    .rt_file_list          (cast_rt_file_list_6_21)
)router_6_21(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_215_to_216),
    .west_valid_i          (valid_215_to_216),
    .west_ready_o          (ready_216_to_215),
    .west_data_o           (data_216_to_215),
    .west_valid_o          (valid_216_to_215),
    .west_ready_i          (ready_215_to_216),
    .east_data_i           (data_217_to_216),
    .east_valid_i          (valid_217_to_216),
    .east_ready_o          (ready_216_to_217),
    .east_data_o           (data_216_to_217),
    .east_valid_o          (valid_216_to_217),
    .east_ready_i          (ready_217_to_216),
    .vert0_data_i          (data_206_to_216_v0),
    .vert0_valid_i         (valid_206_to_216_v0),
    .vert0_ready_o         (ready_216_to_206_v0),
    .vert0_data_o          (data_216_to_226_v0),
    .vert0_valid_o         (valid_216_to_226_v0),
    .vert0_ready_i         (ready_226_to_216_v0),
    .vert1_data_i          (data_206_to_216_v1),
    .vert1_valid_i         (valid_206_to_216_v1),
    .vert1_ready_o         (ready_216_to_206_v1),
    .vert1_data_o          (data_216_to_226_v1),
    .vert1_valid_o         (valid_216_to_226_v1),
    .vert1_ready_i         (ready_226_to_216_v1),
    .local_data_i          (data_i[6][21]),
    .local_valid_i         (valid_i[6][21]),
    .local_ready_o         (ready_o[6][21]),
    .local_data_o          (data_o[6][21]),
    .local_valid_o         (valid_o[6][21]),
    .local_ready_i         (ready_i[6][21]),
    .credit_upd            (credit_upd)
);

/*Router 6,22*/    
cast_router #(
    .isUBM_list            (isUBM_list_6_22),
    .isFC_list             (isFC_list_6_22),
    .FCdn_list             (FCdn_list_6_22),
    .FCpl_list             (FCpl_list_6_22),
    .rt_file_list          (cast_rt_file_list_6_22)
)router_6_22(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_225_to_226),
    .west_valid_i          (valid_225_to_226),
    .west_ready_o          (ready_226_to_225),
    .west_data_o           (data_226_to_225),
    .west_valid_o          (valid_226_to_225),
    .west_ready_i          (ready_225_to_226),
    .east_data_i           (data_227_to_226),
    .east_valid_i          (valid_227_to_226),
    .east_ready_o          (ready_226_to_227),
    .east_data_o           (data_226_to_227),
    .east_valid_o          (valid_226_to_227),
    .east_ready_i          (ready_227_to_226),
    .vert0_data_i          (data_216_to_226_v0),
    .vert0_valid_i         (valid_216_to_226_v0),
    .vert0_ready_o         (ready_226_to_216_v0),
    .vert0_data_o          (data_226_to_236_v0),
    .vert0_valid_o         (valid_226_to_236_v0),
    .vert0_ready_i         (ready_236_to_226_v0),
    .vert1_data_i          (data_216_to_226_v1),
    .vert1_valid_i         (valid_216_to_226_v1),
    .vert1_ready_o         (ready_226_to_216_v1),
    .vert1_data_o          (data_226_to_236_v1),
    .vert1_valid_o         (valid_226_to_236_v1),
    .vert1_ready_i         (ready_236_to_226_v1),
    .local_data_i          (data_i[6][22]),
    .local_valid_i         (valid_i[6][22]),
    .local_ready_o         (ready_o[6][22]),
    .local_data_o          (data_o[6][22]),
    .local_valid_o         (valid_o[6][22]),
    .local_ready_i         (ready_i[6][22]),
    .credit_upd            (credit_upd)
);

/*Router 6,23*/    
cast_router #(
    .isUBM_list            (isUBM_list_6_23),
    .isFC_list             (isFC_list_6_23),
    .FCdn_list             (FCdn_list_6_23),
    .FCpl_list             (FCpl_list_6_23),
    .rt_file_list          (cast_rt_file_list_6_23)
)router_6_23(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_235_to_236),
    .west_valid_i          (valid_235_to_236),
    .west_ready_o          (ready_236_to_235),
    .west_data_o           (data_o_flee3),
    .west_valid_o          (valid_o_flee3),
    .west_ready_i          (ready_i_flee3),
    .east_data_i           (data_237_to_236),
    .east_valid_i          (valid_237_to_236),
    .east_ready_o          (ready_236_to_237),
    .east_data_o           (data_236_to_237),
    .east_valid_o          (valid_236_to_237),
    .east_ready_i          (ready_237_to_236),
    .vert0_data_i          (data_226_to_236_v0),
    .vert0_valid_i         (valid_226_to_236_v0),
    .vert0_ready_o         (ready_236_to_226_v0),
    .vert0_data_o          (data_236_to_246_v0),
    .vert0_valid_o         (valid_236_to_246_v0),
    .vert0_ready_i         (ready_246_to_236_v0),
    .vert1_data_i          (data_226_to_236_v1),
    .vert1_valid_i         (valid_226_to_236_v1),
    .vert1_ready_o         (ready_236_to_226_v1),
    .vert1_data_o          (data_236_to_246_v1),
    .vert1_valid_o         (valid_236_to_246_v1),
    .vert1_ready_i         (ready_246_to_236_v1),
    .local_data_i          (data_i[6][23]),
    .local_valid_i         (valid_i[6][23]),
    .local_ready_o         (ready_o[6][23]),
    .local_data_o          (data_o[6][23]),
    .local_valid_o         (valid_o[6][23]),
    .local_ready_i         (ready_i[6][23]),
    .credit_upd            (credit_upd)
);

/*Router 6,24*/    
cast_router #(
    .isUBM_list            (isUBM_list_6_24),
    .isFC_list             (isFC_list_6_24),
    .FCdn_list             (FCdn_list_6_24),
    .FCpl_list             (FCpl_list_6_24),
    .rt_file_list          (cast_rt_file_list_6_24)
)router_6_24(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_245_to_246),
    .west_valid_i          (valid_245_to_246),
    .west_ready_o          (ready_246_to_245),
    .west_data_o           (data_246_to_245),
    .west_valid_o          (valid_246_to_245),
    .west_ready_i          (ready_245_to_246),
    .east_data_i           (data_247_to_246),
    .east_valid_i          (valid_247_to_246),
    .east_ready_o          (ready_246_to_247),
    .east_data_o           (data_246_to_247),
    .east_valid_o          (valid_246_to_247),
    .east_ready_i          (ready_247_to_246),
    .vert0_data_i          (data_236_to_246_v0),
    .vert0_valid_i         (valid_236_to_246_v0),
    .vert0_ready_o         (ready_246_to_236_v0),
    .vert0_data_o          (),
    .vert0_valid_o         (),
    .vert0_ready_i         (1'b0),
    .vert1_data_i          (data_236_to_246_v1),
    .vert1_valid_i         (valid_236_to_246_v1),
    .vert1_ready_o         (ready_246_to_236_v1),
    .vert1_data_o          (),
    .vert1_valid_o         (),
    .vert1_ready_i         (1'b0),
    .local_data_i          (data_i[6][24]),
    .local_valid_i         (valid_i[6][24]),
    .local_ready_o         (ready_o[6][24]),
    .local_data_o          (data_o[6][24]),
    .local_valid_o         (valid_o[6][24]),
    .local_ready_i         (ready_i[6][24]),
    .credit_upd            (credit_upd)
);

/*Router 7,0*/    
cast_router #(
    .isUBM_list            (isUBM_list_7_0),
    .isFC_list             (isFC_list_7_0),
    .FCdn_list             (FCdn_list_7_0),
    .FCpl_list             (FCpl_list_7_0),
    .rt_file_list          (cast_rt_file_list_7_0)
)router_7_0(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_6_to_7),
    .west_valid_i          (valid_6_to_7),
    .west_ready_o          (ready_7_to_6),
    .west_data_o           (data_7_to_6),
    .west_valid_o          (valid_7_to_6),
    .west_ready_i          (ready_6_to_7),
    .east_data_i           (data_8_to_7),
    .east_valid_i          (valid_8_to_7),
    .east_ready_o          (ready_7_to_8),
    .east_data_o           (data_7_to_8),
    .east_valid_o          (valid_7_to_8),
    .east_ready_i          (ready_8_to_7),
    .vert0_data_i          (34'b0),
    .vert0_valid_i         (1'b0),
    .vert0_ready_o         (),
    .vert0_data_o          (data_7_to_17_v0),
    .vert0_valid_o         (valid_7_to_17_v0),
    .vert0_ready_i         (ready_17_to_7_v0),
    .vert1_data_i          (34'b0),
    .vert1_valid_i         (1'b0),
    .vert1_ready_o         (),
    .vert1_data_o          (data_7_to_17_v1),
    .vert1_valid_o         (valid_7_to_17_v1),
    .vert1_ready_i         (ready_17_to_7_v1),
    .local_data_i          (data_i[7][0]),
    .local_valid_i         (valid_i[7][0]),
    .local_ready_o         (ready_o[7][0]),
    .local_data_o          (data_o[7][0]),
    .local_valid_o         (valid_o[7][0]),
    .local_ready_i         (ready_i[7][0]),
    .credit_upd            (credit_upd)
);

/*Router 7,1*/    
cast_router #(
    .isUBM_list            (isUBM_list_7_1),
    .isFC_list             (isFC_list_7_1),
    .FCdn_list             (FCdn_list_7_1),
    .FCpl_list             (FCpl_list_7_1),
    .rt_file_list          (cast_rt_file_list_7_1)
)router_7_1(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_16_to_17),
    .west_valid_i          (valid_16_to_17),
    .west_ready_o          (ready_17_to_16),
    .west_data_o           (data_17_to_16),
    .west_valid_o          (valid_17_to_16),
    .west_ready_i          (ready_16_to_17),
    .east_data_i           (data_18_to_17),
    .east_valid_i          (valid_18_to_17),
    .east_ready_o          (ready_17_to_18),
    .east_data_o           (data_17_to_18),
    .east_valid_o          (valid_17_to_18),
    .east_ready_i          (ready_18_to_17),
    .vert0_data_i          (data_7_to_17_v0),
    .vert0_valid_i         (valid_7_to_17_v0),
    .vert0_ready_o         (ready_17_to_7_v0),
    .vert0_data_o          (data_17_to_27_v0),
    .vert0_valid_o         (valid_17_to_27_v0),
    .vert0_ready_i         (ready_27_to_17_v0),
    .vert1_data_i          (data_7_to_17_v1),
    .vert1_valid_i         (valid_7_to_17_v1),
    .vert1_ready_o         (ready_17_to_7_v1),
    .vert1_data_o          (data_17_to_27_v1),
    .vert1_valid_o         (valid_17_to_27_v1),
    .vert1_ready_i         (ready_27_to_17_v1),
    .local_data_i          (data_i[7][1]),
    .local_valid_i         (valid_i[7][1]),
    .local_ready_o         (ready_o[7][1]),
    .local_data_o          (data_o[7][1]),
    .local_valid_o         (valid_o[7][1]),
    .local_ready_i         (ready_i[7][1]),
    .credit_upd            (credit_upd)
);

/*Router 7,2*/    
cast_router #(
    .isUBM_list            (isUBM_list_7_2),
    .isFC_list             (isFC_list_7_2),
    .FCdn_list             (FCdn_list_7_2),
    .FCpl_list             (FCpl_list_7_2),
    .rt_file_list          (cast_rt_file_list_7_2)
)router_7_2(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_26_to_27),
    .west_valid_i          (valid_26_to_27),
    .west_ready_o          (ready_27_to_26),
    .west_data_o           (data_27_to_26),
    .west_valid_o          (valid_27_to_26),
    .west_ready_i          (ready_26_to_27),
    .east_data_i           (data_28_to_27),
    .east_valid_i          (valid_28_to_27),
    .east_ready_o          (ready_27_to_28),
    .east_data_o           (data_27_to_28),
    .east_valid_o          (valid_27_to_28),
    .east_ready_i          (ready_28_to_27),
    .vert0_data_i          (data_17_to_27_v0),
    .vert0_valid_i         (valid_17_to_27_v0),
    .vert0_ready_o         (ready_27_to_17_v0),
    .vert0_data_o          (data_27_to_37_v0),
    .vert0_valid_o         (valid_27_to_37_v0),
    .vert0_ready_i         (ready_37_to_27_v0),
    .vert1_data_i          (data_17_to_27_v1),
    .vert1_valid_i         (valid_17_to_27_v1),
    .vert1_ready_o         (ready_27_to_17_v1),
    .vert1_data_o          (data_27_to_37_v1),
    .vert1_valid_o         (valid_27_to_37_v1),
    .vert1_ready_i         (ready_37_to_27_v1),
    .local_data_i          (data_i[7][2]),
    .local_valid_i         (valid_i[7][2]),
    .local_ready_o         (ready_o[7][2]),
    .local_data_o          (data_o[7][2]),
    .local_valid_o         (valid_o[7][2]),
    .local_ready_i         (ready_i[7][2]),
    .credit_upd            (credit_upd)
);

/*Router 7,3*/    
cast_router #(
    .isUBM_list            (isUBM_list_7_3),
    .isFC_list             (isFC_list_7_3),
    .FCdn_list             (FCdn_list_7_3),
    .FCpl_list             (FCpl_list_7_3),
    .rt_file_list          (cast_rt_file_list_7_3)
)router_7_3(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_36_to_37),
    .west_valid_i          (valid_36_to_37),
    .west_ready_o          (ready_37_to_36),
    .west_data_o           (data_37_to_36),
    .west_valid_o          (valid_37_to_36),
    .west_ready_i          (ready_36_to_37),
    .east_data_i           (data_38_to_37),
    .east_valid_i          (valid_38_to_37),
    .east_ready_o          (ready_37_to_38),
    .east_data_o           (data_37_to_38),
    .east_valid_o          (valid_37_to_38),
    .east_ready_i          (ready_38_to_37),
    .vert0_data_i          (data_27_to_37_v0),
    .vert0_valid_i         (valid_27_to_37_v0),
    .vert0_ready_o         (ready_37_to_27_v0),
    .vert0_data_o          (data_37_to_47_v0),
    .vert0_valid_o         (valid_37_to_47_v0),
    .vert0_ready_i         (ready_47_to_37_v0),
    .vert1_data_i          (data_27_to_37_v1),
    .vert1_valid_i         (valid_27_to_37_v1),
    .vert1_ready_o         (ready_37_to_27_v1),
    .vert1_data_o          (data_37_to_47_v1),
    .vert1_valid_o         (valid_37_to_47_v1),
    .vert1_ready_i         (ready_47_to_37_v1),
    .local_data_i          (data_i[7][3]),
    .local_valid_i         (valid_i[7][3]),
    .local_ready_o         (ready_o[7][3]),
    .local_data_o          (data_o[7][3]),
    .local_valid_o         (valid_o[7][3]),
    .local_ready_i         (ready_i[7][3]),
    .credit_upd            (credit_upd)
);

/*Router 7,4*/    
cast_router #(
    .isUBM_list            (isUBM_list_7_4),
    .isFC_list             (isFC_list_7_4),
    .FCdn_list             (FCdn_list_7_4),
    .FCpl_list             (FCpl_list_7_4),
    .rt_file_list          (cast_rt_file_list_7_4)
)router_7_4(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_46_to_47),
    .west_valid_i          (valid_46_to_47),
    .west_ready_o          (ready_47_to_46),
    .west_data_o           (data_47_to_46),
    .west_valid_o          (valid_47_to_46),
    .west_ready_i          (ready_46_to_47),
    .east_data_i           (data_48_to_47),
    .east_valid_i          (valid_48_to_47),
    .east_ready_o          (ready_47_to_48),
    .east_data_o           (data_47_to_48),
    .east_valid_o          (valid_47_to_48),
    .east_ready_i          (ready_48_to_47),
    .vert0_data_i          (data_37_to_47_v0),
    .vert0_valid_i         (valid_37_to_47_v0),
    .vert0_ready_o         (ready_47_to_37_v0),
    .vert0_data_o          (data_47_to_57_v0),
    .vert0_valid_o         (valid_47_to_57_v0),
    .vert0_ready_i         (ready_57_to_47_v0),
    .vert1_data_i          (data_37_to_47_v1),
    .vert1_valid_i         (valid_37_to_47_v1),
    .vert1_ready_o         (ready_47_to_37_v1),
    .vert1_data_o          (data_47_to_57_v1),
    .vert1_valid_o         (valid_47_to_57_v1),
    .vert1_ready_i         (ready_57_to_47_v1),
    .local_data_i          (data_i[7][4]),
    .local_valid_i         (valid_i[7][4]),
    .local_ready_o         (ready_o[7][4]),
    .local_data_o          (data_o[7][4]),
    .local_valid_o         (valid_o[7][4]),
    .local_ready_i         (ready_i[7][4]),
    .credit_upd            (credit_upd)
);

/*Router 7,5*/    
cast_router #(
    .isUBM_list            (isUBM_list_7_5),
    .isFC_list             (isFC_list_7_5),
    .FCdn_list             (FCdn_list_7_5),
    .FCpl_list             (FCpl_list_7_5),
    .rt_file_list          (cast_rt_file_list_7_5)
)router_7_5(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_56_to_57),
    .west_valid_i          (valid_56_to_57),
    .west_ready_o          (ready_57_to_56),
    .west_data_o           (data_57_to_56),
    .west_valid_o          (valid_57_to_56),
    .west_ready_i          (ready_56_to_57),
    .east_data_i           (data_58_to_57),
    .east_valid_i          (valid_58_to_57),
    .east_ready_o          (ready_57_to_58),
    .east_data_o           (data_57_to_58),
    .east_valid_o          (valid_57_to_58),
    .east_ready_i          (ready_58_to_57),
    .vert0_data_i          (data_47_to_57_v0),
    .vert0_valid_i         (valid_47_to_57_v0),
    .vert0_ready_o         (ready_57_to_47_v0),
    .vert0_data_o          (data_57_to_67_v0),
    .vert0_valid_o         (valid_57_to_67_v0),
    .vert0_ready_i         (ready_67_to_57_v0),
    .vert1_data_i          (data_47_to_57_v1),
    .vert1_valid_i         (valid_47_to_57_v1),
    .vert1_ready_o         (ready_57_to_47_v1),
    .vert1_data_o          (data_57_to_67_v1),
    .vert1_valid_o         (valid_57_to_67_v1),
    .vert1_ready_i         (ready_67_to_57_v1),
    .local_data_i          (data_i[7][5]),
    .local_valid_i         (valid_i[7][5]),
    .local_ready_o         (ready_o[7][5]),
    .local_data_o          (data_o[7][5]),
    .local_valid_o         (valid_o[7][5]),
    .local_ready_i         (ready_i[7][5]),
    .credit_upd            (credit_upd)
);

/*Router 7,6*/    
cast_router #(
    .isUBM_list            (isUBM_list_7_6),
    .isFC_list             (isFC_list_7_6),
    .FCdn_list             (FCdn_list_7_6),
    .FCpl_list             (FCpl_list_7_6),
    .rt_file_list          (cast_rt_file_list_7_6)
)router_7_6(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_66_to_67),
    .west_valid_i          (valid_66_to_67),
    .west_ready_o          (ready_67_to_66),
    .west_data_o           (data_67_to_66),
    .west_valid_o          (valid_67_to_66),
    .west_ready_i          (ready_66_to_67),
    .east_data_i           (data_68_to_67),
    .east_valid_i          (valid_68_to_67),
    .east_ready_o          (ready_67_to_68),
    .east_data_o           (data_67_to_68),
    .east_valid_o          (valid_67_to_68),
    .east_ready_i          (ready_68_to_67),
    .vert0_data_i          (data_57_to_67_v0),
    .vert0_valid_i         (valid_57_to_67_v0),
    .vert0_ready_o         (ready_67_to_57_v0),
    .vert0_data_o          (data_67_to_77_v0),
    .vert0_valid_o         (valid_67_to_77_v0),
    .vert0_ready_i         (ready_77_to_67_v0),
    .vert1_data_i          (data_57_to_67_v1),
    .vert1_valid_i         (valid_57_to_67_v1),
    .vert1_ready_o         (ready_67_to_57_v1),
    .vert1_data_o          (data_67_to_77_v1),
    .vert1_valid_o         (valid_67_to_77_v1),
    .vert1_ready_i         (ready_77_to_67_v1),
    .local_data_i          (data_i[7][6]),
    .local_valid_i         (valid_i[7][6]),
    .local_ready_o         (ready_o[7][6]),
    .local_data_o          (data_o[7][6]),
    .local_valid_o         (valid_o[7][6]),
    .local_ready_i         (ready_i[7][6]),
    .credit_upd            (credit_upd)
);

/*Router 7,7*/    
cast_router #(
    .isUBM_list            (isUBM_list_7_7),
    .isFC_list             (isFC_list_7_7),
    .FCdn_list             (FCdn_list_7_7),
    .FCpl_list             (FCpl_list_7_7),
    .rt_file_list          (cast_rt_file_list_7_7)
)router_7_7(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_76_to_77),
    .west_valid_i          (valid_76_to_77),
    .west_ready_o          (ready_77_to_76),
    .west_data_o           (data_77_to_76),
    .west_valid_o          (valid_77_to_76),
    .west_ready_i          (ready_76_to_77),
    .east_data_i           (data_78_to_77),
    .east_valid_i          (valid_78_to_77),
    .east_ready_o          (ready_77_to_78),
    .east_data_o           (data_77_to_78),
    .east_valid_o          (valid_77_to_78),
    .east_ready_i          (ready_78_to_77),
    .vert0_data_i          (data_67_to_77_v0),
    .vert0_valid_i         (valid_67_to_77_v0),
    .vert0_ready_o         (ready_77_to_67_v0),
    .vert0_data_o          (data_77_to_87_v0),
    .vert0_valid_o         (valid_77_to_87_v0),
    .vert0_ready_i         (ready_87_to_77_v0),
    .vert1_data_i          (data_67_to_77_v1),
    .vert1_valid_i         (valid_67_to_77_v1),
    .vert1_ready_o         (ready_77_to_67_v1),
    .vert1_data_o          (data_77_to_87_v1),
    .vert1_valid_o         (valid_77_to_87_v1),
    .vert1_ready_i         (ready_87_to_77_v1),
    .local_data_i          (data_i[7][7]),
    .local_valid_i         (valid_i[7][7]),
    .local_ready_o         (ready_o[7][7]),
    .local_data_o          (data_o[7][7]),
    .local_valid_o         (valid_o[7][7]),
    .local_ready_i         (ready_i[7][7]),
    .credit_upd            (credit_upd)
);

/*Router 7,8*/    
cast_router #(
    .isUBM_list            (isUBM_list_7_8),
    .isFC_list             (isFC_list_7_8),
    .FCdn_list             (FCdn_list_7_8),
    .FCpl_list             (FCpl_list_7_8),
    .rt_file_list          (cast_rt_file_list_7_8)
)router_7_8(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_86_to_87),
    .west_valid_i          (valid_86_to_87),
    .west_ready_o          (ready_87_to_86),
    .west_data_o           (data_87_to_86),
    .west_valid_o          (valid_87_to_86),
    .west_ready_i          (ready_86_to_87),
    .east_data_i           (data_88_to_87),
    .east_valid_i          (valid_88_to_87),
    .east_ready_o          (ready_87_to_88),
    .east_data_o           (data_87_to_88),
    .east_valid_o          (valid_87_to_88),
    .east_ready_i          (ready_88_to_87),
    .vert0_data_i          (data_77_to_87_v0),
    .vert0_valid_i         (valid_77_to_87_v0),
    .vert0_ready_o         (ready_87_to_77_v0),
    .vert0_data_o          (data_87_to_97_v0),
    .vert0_valid_o         (valid_87_to_97_v0),
    .vert0_ready_i         (ready_97_to_87_v0),
    .vert1_data_i          (data_77_to_87_v1),
    .vert1_valid_i         (valid_77_to_87_v1),
    .vert1_ready_o         (ready_87_to_77_v1),
    .vert1_data_o          (data_87_to_97_v1),
    .vert1_valid_o         (valid_87_to_97_v1),
    .vert1_ready_i         (ready_97_to_87_v1),
    .local_data_i          (data_i[7][8]),
    .local_valid_i         (valid_i[7][8]),
    .local_ready_o         (ready_o[7][8]),
    .local_data_o          (data_o[7][8]),
    .local_valid_o         (valid_o[7][8]),
    .local_ready_i         (ready_i[7][8]),
    .credit_upd            (credit_upd)
);

/*Router 7,9*/    
cast_router #(
    .isUBM_list            (isUBM_list_7_9),
    .isFC_list             (isFC_list_7_9),
    .FCdn_list             (FCdn_list_7_9),
    .FCpl_list             (FCpl_list_7_9),
    .rt_file_list          (cast_rt_file_list_7_9)
)router_7_9(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_96_to_97),
    .west_valid_i          (valid_96_to_97),
    .west_ready_o          (ready_97_to_96),
    .west_data_o           (data_97_to_96),
    .west_valid_o          (valid_97_to_96),
    .west_ready_i          (ready_96_to_97),
    .east_data_i           (data_98_to_97),
    .east_valid_i          (valid_98_to_97),
    .east_ready_o          (ready_97_to_98),
    .east_data_o           (data_97_to_98),
    .east_valid_o          (valid_97_to_98),
    .east_ready_i          (ready_98_to_97),
    .vert0_data_i          (data_87_to_97_v0),
    .vert0_valid_i         (valid_87_to_97_v0),
    .vert0_ready_o         (ready_97_to_87_v0),
    .vert0_data_o          (data_97_to_107_v0),
    .vert0_valid_o         (valid_97_to_107_v0),
    .vert0_ready_i         (ready_107_to_97_v0),
    .vert1_data_i          (data_87_to_97_v1),
    .vert1_valid_i         (valid_87_to_97_v1),
    .vert1_ready_o         (ready_97_to_87_v1),
    .vert1_data_o          (data_97_to_107_v1),
    .vert1_valid_o         (valid_97_to_107_v1),
    .vert1_ready_i         (ready_107_to_97_v1),
    .local_data_i          (data_i[7][9]),
    .local_valid_i         (valid_i[7][9]),
    .local_ready_o         (ready_o[7][9]),
    .local_data_o          (data_o[7][9]),
    .local_valid_o         (valid_o[7][9]),
    .local_ready_i         (ready_i[7][9]),
    .credit_upd            (credit_upd)
);

/*Router 7,10*/    
cast_router #(
    .isUBM_list            (isUBM_list_7_10),
    .isFC_list             (isFC_list_7_10),
    .FCdn_list             (FCdn_list_7_10),
    .FCpl_list             (FCpl_list_7_10),
    .rt_file_list          (cast_rt_file_list_7_10)
)router_7_10(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_106_to_107),
    .west_valid_i          (valid_106_to_107),
    .west_ready_o          (ready_107_to_106),
    .west_data_o           (data_107_to_106),
    .west_valid_o          (valid_107_to_106),
    .west_ready_i          (ready_106_to_107),
    .east_data_i           (data_108_to_107),
    .east_valid_i          (valid_108_to_107),
    .east_ready_o          (ready_107_to_108),
    .east_data_o           (data_107_to_108),
    .east_valid_o          (valid_107_to_108),
    .east_ready_i          (ready_108_to_107),
    .vert0_data_i          (data_97_to_107_v0),
    .vert0_valid_i         (valid_97_to_107_v0),
    .vert0_ready_o         (ready_107_to_97_v0),
    .vert0_data_o          (data_107_to_117_v0),
    .vert0_valid_o         (valid_107_to_117_v0),
    .vert0_ready_i         (ready_117_to_107_v0),
    .vert1_data_i          (data_97_to_107_v1),
    .vert1_valid_i         (valid_97_to_107_v1),
    .vert1_ready_o         (ready_107_to_97_v1),
    .vert1_data_o          (data_107_to_117_v1),
    .vert1_valid_o         (valid_107_to_117_v1),
    .vert1_ready_i         (ready_117_to_107_v1),
    .local_data_i          (data_i[7][10]),
    .local_valid_i         (valid_i[7][10]),
    .local_ready_o         (ready_o[7][10]),
    .local_data_o          (data_o[7][10]),
    .local_valid_o         (valid_o[7][10]),
    .local_ready_i         (ready_i[7][10]),
    .credit_upd            (credit_upd)
);

/*Router 7,11*/    
cast_router #(
    .isUBM_list            (isUBM_list_7_11),
    .isFC_list             (isFC_list_7_11),
    .FCdn_list             (FCdn_list_7_11),
    .FCpl_list             (FCpl_list_7_11),
    .rt_file_list          (cast_rt_file_list_7_11)
)router_7_11(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_116_to_117),
    .west_valid_i          (valid_116_to_117),
    .west_ready_o          (ready_117_to_116),
    .west_data_o           (data_117_to_116),
    .west_valid_o          (valid_117_to_116),
    .west_ready_i          (ready_116_to_117),
    .east_data_i           (data_118_to_117),
    .east_valid_i          (valid_118_to_117),
    .east_ready_o          (ready_117_to_118),
    .east_data_o           (data_117_to_118),
    .east_valid_o          (valid_117_to_118),
    .east_ready_i          (ready_118_to_117),
    .vert0_data_i          (data_107_to_117_v0),
    .vert0_valid_i         (valid_107_to_117_v0),
    .vert0_ready_o         (ready_117_to_107_v0),
    .vert0_data_o          (data_117_to_127_v0),
    .vert0_valid_o         (valid_117_to_127_v0),
    .vert0_ready_i         (ready_127_to_117_v0),
    .vert1_data_i          (data_107_to_117_v1),
    .vert1_valid_i         (valid_107_to_117_v1),
    .vert1_ready_o         (ready_117_to_107_v1),
    .vert1_data_o          (data_117_to_127_v1),
    .vert1_valid_o         (valid_117_to_127_v1),
    .vert1_ready_i         (ready_127_to_117_v1),
    .local_data_i          (data_i[7][11]),
    .local_valid_i         (valid_i[7][11]),
    .local_ready_o         (ready_o[7][11]),
    .local_data_o          (data_o[7][11]),
    .local_valid_o         (valid_o[7][11]),
    .local_ready_i         (ready_i[7][11]),
    .credit_upd            (credit_upd)
);

/*Router 7,12*/    
cast_router #(
    .isUBM_list            (isUBM_list_7_12),
    .isFC_list             (isFC_list_7_12),
    .FCdn_list             (FCdn_list_7_12),
    .FCpl_list             (FCpl_list_7_12),
    .rt_file_list          (cast_rt_file_list_7_12)
)router_7_12(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_126_to_127),
    .west_valid_i          (valid_126_to_127),
    .west_ready_o          (ready_127_to_126),
    .west_data_o           (data_127_to_126),
    .west_valid_o          (valid_127_to_126),
    .west_ready_i          (ready_126_to_127),
    .east_data_i           (data_128_to_127),
    .east_valid_i          (valid_128_to_127),
    .east_ready_o          (ready_127_to_128),
    .east_data_o           (data_127_to_128),
    .east_valid_o          (valid_127_to_128),
    .east_ready_i          (ready_128_to_127),
    .vert0_data_i          (data_117_to_127_v0),
    .vert0_valid_i         (valid_117_to_127_v0),
    .vert0_ready_o         (ready_127_to_117_v0),
    .vert0_data_o          (data_127_to_137_v0),
    .vert0_valid_o         (valid_127_to_137_v0),
    .vert0_ready_i         (ready_137_to_127_v0),
    .vert1_data_i          (data_117_to_127_v1),
    .vert1_valid_i         (valid_117_to_127_v1),
    .vert1_ready_o         (ready_127_to_117_v1),
    .vert1_data_o          (data_127_to_137_v1),
    .vert1_valid_o         (valid_127_to_137_v1),
    .vert1_ready_i         (ready_137_to_127_v1),
    .local_data_i          (data_i[7][12]),
    .local_valid_i         (valid_i[7][12]),
    .local_ready_o         (ready_o[7][12]),
    .local_data_o          (data_o[7][12]),
    .local_valid_o         (valid_o[7][12]),
    .local_ready_i         (ready_i[7][12]),
    .credit_upd            (credit_upd)
);

/*Router 7,13*/    
cast_router #(
    .isUBM_list            (isUBM_list_7_13),
    .isFC_list             (isFC_list_7_13),
    .FCdn_list             (FCdn_list_7_13),
    .FCpl_list             (FCpl_list_7_13),
    .rt_file_list          (cast_rt_file_list_7_13)
)router_7_13(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_136_to_137),
    .west_valid_i          (valid_136_to_137),
    .west_ready_o          (ready_137_to_136),
    .west_data_o           (data_137_to_136),
    .west_valid_o          (valid_137_to_136),
    .west_ready_i          (ready_136_to_137),
    .east_data_i           (data_138_to_137),
    .east_valid_i          (valid_138_to_137),
    .east_ready_o          (ready_137_to_138),
    .east_data_o           (data_137_to_138),
    .east_valid_o          (valid_137_to_138),
    .east_ready_i          (ready_138_to_137),
    .vert0_data_i          (data_127_to_137_v0),
    .vert0_valid_i         (valid_127_to_137_v0),
    .vert0_ready_o         (ready_137_to_127_v0),
    .vert0_data_o          (data_137_to_147_v0),
    .vert0_valid_o         (valid_137_to_147_v0),
    .vert0_ready_i         (ready_147_to_137_v0),
    .vert1_data_i          (data_127_to_137_v1),
    .vert1_valid_i         (valid_127_to_137_v1),
    .vert1_ready_o         (ready_137_to_127_v1),
    .vert1_data_o          (data_137_to_147_v1),
    .vert1_valid_o         (valid_137_to_147_v1),
    .vert1_ready_i         (ready_147_to_137_v1),
    .local_data_i          (data_i[7][13]),
    .local_valid_i         (valid_i[7][13]),
    .local_ready_o         (ready_o[7][13]),
    .local_data_o          (data_o[7][13]),
    .local_valid_o         (valid_o[7][13]),
    .local_ready_i         (ready_i[7][13]),
    .credit_upd            (credit_upd)
);

/*Router 7,14*/    
cast_router #(
    .isUBM_list            (isUBM_list_7_14),
    .isFC_list             (isFC_list_7_14),
    .FCdn_list             (FCdn_list_7_14),
    .FCpl_list             (FCpl_list_7_14),
    .rt_file_list          (cast_rt_file_list_7_14)
)router_7_14(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_146_to_147),
    .west_valid_i          (valid_146_to_147),
    .west_ready_o          (ready_147_to_146),
    .west_data_o           (data_147_to_146),
    .west_valid_o          (valid_147_to_146),
    .west_ready_i          (ready_146_to_147),
    .east_data_i           (data_148_to_147),
    .east_valid_i          (valid_148_to_147),
    .east_ready_o          (ready_147_to_148),
    .east_data_o           (data_147_to_148),
    .east_valid_o          (valid_147_to_148),
    .east_ready_i          (ready_148_to_147),
    .vert0_data_i          (data_137_to_147_v0),
    .vert0_valid_i         (valid_137_to_147_v0),
    .vert0_ready_o         (ready_147_to_137_v0),
    .vert0_data_o          (data_147_to_157_v0),
    .vert0_valid_o         (valid_147_to_157_v0),
    .vert0_ready_i         (ready_157_to_147_v0),
    .vert1_data_i          (data_137_to_147_v1),
    .vert1_valid_i         (valid_137_to_147_v1),
    .vert1_ready_o         (ready_147_to_137_v1),
    .vert1_data_o          (data_147_to_157_v1),
    .vert1_valid_o         (valid_147_to_157_v1),
    .vert1_ready_i         (ready_157_to_147_v1),
    .local_data_i          (data_i[7][14]),
    .local_valid_i         (valid_i[7][14]),
    .local_ready_o         (ready_o[7][14]),
    .local_data_o          (data_o[7][14]),
    .local_valid_o         (valid_o[7][14]),
    .local_ready_i         (ready_i[7][14]),
    .credit_upd            (credit_upd)
);

/*Router 7,15*/    
cast_router #(
    .isUBM_list            (isUBM_list_7_15),
    .isFC_list             (isFC_list_7_15),
    .FCdn_list             (FCdn_list_7_15),
    .FCpl_list             (FCpl_list_7_15),
    .rt_file_list          (cast_rt_file_list_7_15)
)router_7_15(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_156_to_157),
    .west_valid_i          (valid_156_to_157),
    .west_ready_o          (ready_157_to_156),
    .west_data_o           (data_157_to_156),
    .west_valid_o          (valid_157_to_156),
    .west_ready_i          (ready_156_to_157),
    .east_data_i           (data_158_to_157),
    .east_valid_i          (valid_158_to_157),
    .east_ready_o          (ready_157_to_158),
    .east_data_o           (data_157_to_158),
    .east_valid_o          (valid_157_to_158),
    .east_ready_i          (ready_158_to_157),
    .vert0_data_i          (data_147_to_157_v0),
    .vert0_valid_i         (valid_147_to_157_v0),
    .vert0_ready_o         (ready_157_to_147_v0),
    .vert0_data_o          (data_157_to_167_v0),
    .vert0_valid_o         (valid_157_to_167_v0),
    .vert0_ready_i         (ready_167_to_157_v0),
    .vert1_data_i          (data_147_to_157_v1),
    .vert1_valid_i         (valid_147_to_157_v1),
    .vert1_ready_o         (ready_157_to_147_v1),
    .vert1_data_o          (data_157_to_167_v1),
    .vert1_valid_o         (valid_157_to_167_v1),
    .vert1_ready_i         (ready_167_to_157_v1),
    .local_data_i          (data_i[7][15]),
    .local_valid_i         (valid_i[7][15]),
    .local_ready_o         (ready_o[7][15]),
    .local_data_o          (data_o[7][15]),
    .local_valid_o         (valid_o[7][15]),
    .local_ready_i         (ready_i[7][15]),
    .credit_upd            (credit_upd)
);

/*Router 7,16*/    
cast_router #(
    .isUBM_list            (isUBM_list_7_16),
    .isFC_list             (isFC_list_7_16),
    .FCdn_list             (FCdn_list_7_16),
    .FCpl_list             (FCpl_list_7_16),
    .rt_file_list          (cast_rt_file_list_7_16)
)router_7_16(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_166_to_167),
    .west_valid_i          (valid_166_to_167),
    .west_ready_o          (ready_167_to_166),
    .west_data_o           (data_167_to_166),
    .west_valid_o          (valid_167_to_166),
    .west_ready_i          (ready_166_to_167),
    .east_data_i           (data_168_to_167),
    .east_valid_i          (valid_168_to_167),
    .east_ready_o          (ready_167_to_168),
    .east_data_o           (data_167_to_168),
    .east_valid_o          (valid_167_to_168),
    .east_ready_i          (ready_168_to_167),
    .vert0_data_i          (data_157_to_167_v0),
    .vert0_valid_i         (valid_157_to_167_v0),
    .vert0_ready_o         (ready_167_to_157_v0),
    .vert0_data_o          (data_167_to_177_v0),
    .vert0_valid_o         (valid_167_to_177_v0),
    .vert0_ready_i         (ready_177_to_167_v0),
    .vert1_data_i          (data_157_to_167_v1),
    .vert1_valid_i         (valid_157_to_167_v1),
    .vert1_ready_o         (ready_167_to_157_v1),
    .vert1_data_o          (data_167_to_177_v1),
    .vert1_valid_o         (valid_167_to_177_v1),
    .vert1_ready_i         (ready_177_to_167_v1),
    .local_data_i          (data_i[7][16]),
    .local_valid_i         (valid_i[7][16]),
    .local_ready_o         (ready_o[7][16]),
    .local_data_o          (data_o[7][16]),
    .local_valid_o         (valid_o[7][16]),
    .local_ready_i         (ready_i[7][16]),
    .credit_upd            (credit_upd)
);

/*Router 7,17*/    
cast_router #(
    .isUBM_list            (isUBM_list_7_17),
    .isFC_list             (isFC_list_7_17),
    .FCdn_list             (FCdn_list_7_17),
    .FCpl_list             (FCpl_list_7_17),
    .rt_file_list          (cast_rt_file_list_7_17)
)router_7_17(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_176_to_177),
    .west_valid_i          (valid_176_to_177),
    .west_ready_o          (ready_177_to_176),
    .west_data_o           (data_177_to_176),
    .west_valid_o          (valid_177_to_176),
    .west_ready_i          (ready_176_to_177),
    .east_data_i           (data_178_to_177),
    .east_valid_i          (valid_178_to_177),
    .east_ready_o          (ready_177_to_178),
    .east_data_o           (data_177_to_178),
    .east_valid_o          (valid_177_to_178),
    .east_ready_i          (ready_178_to_177),
    .vert0_data_i          (data_167_to_177_v0),
    .vert0_valid_i         (valid_167_to_177_v0),
    .vert0_ready_o         (ready_177_to_167_v0),
    .vert0_data_o          (data_177_to_187_v0),
    .vert0_valid_o         (valid_177_to_187_v0),
    .vert0_ready_i         (ready_187_to_177_v0),
    .vert1_data_i          (data_167_to_177_v1),
    .vert1_valid_i         (valid_167_to_177_v1),
    .vert1_ready_o         (ready_177_to_167_v1),
    .vert1_data_o          (data_177_to_187_v1),
    .vert1_valid_o         (valid_177_to_187_v1),
    .vert1_ready_i         (ready_187_to_177_v1),
    .local_data_i          (data_i[7][17]),
    .local_valid_i         (valid_i[7][17]),
    .local_ready_o         (ready_o[7][17]),
    .local_data_o          (data_o[7][17]),
    .local_valid_o         (valid_o[7][17]),
    .local_ready_i         (ready_i[7][17]),
    .credit_upd            (credit_upd)
);

/*Router 7,18*/    
cast_router #(
    .isUBM_list            (isUBM_list_7_18),
    .isFC_list             (isFC_list_7_18),
    .FCdn_list             (FCdn_list_7_18),
    .FCpl_list             (FCpl_list_7_18),
    .rt_file_list          (cast_rt_file_list_7_18)
)router_7_18(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_186_to_187),
    .west_valid_i          (valid_186_to_187),
    .west_ready_o          (ready_187_to_186),
    .west_data_o           (data_187_to_186),
    .west_valid_o          (valid_187_to_186),
    .west_ready_i          (ready_186_to_187),
    .east_data_i           (data_188_to_187),
    .east_valid_i          (valid_188_to_187),
    .east_ready_o          (ready_187_to_188),
    .east_data_o           (data_187_to_188),
    .east_valid_o          (valid_187_to_188),
    .east_ready_i          (ready_188_to_187),
    .vert0_data_i          (data_177_to_187_v0),
    .vert0_valid_i         (valid_177_to_187_v0),
    .vert0_ready_o         (ready_187_to_177_v0),
    .vert0_data_o          (data_187_to_197_v0),
    .vert0_valid_o         (valid_187_to_197_v0),
    .vert0_ready_i         (ready_197_to_187_v0),
    .vert1_data_i          (data_177_to_187_v1),
    .vert1_valid_i         (valid_177_to_187_v1),
    .vert1_ready_o         (ready_187_to_177_v1),
    .vert1_data_o          (data_187_to_197_v1),
    .vert1_valid_o         (valid_187_to_197_v1),
    .vert1_ready_i         (ready_197_to_187_v1),
    .local_data_i          (data_i[7][18]),
    .local_valid_i         (valid_i[7][18]),
    .local_ready_o         (ready_o[7][18]),
    .local_data_o          (data_o[7][18]),
    .local_valid_o         (valid_o[7][18]),
    .local_ready_i         (ready_i[7][18]),
    .credit_upd            (credit_upd)
);

/*Router 7,19*/    
cast_router #(
    .isUBM_list            (isUBM_list_7_19),
    .isFC_list             (isFC_list_7_19),
    .FCdn_list             (FCdn_list_7_19),
    .FCpl_list             (FCpl_list_7_19),
    .rt_file_list          (cast_rt_file_list_7_19)
)router_7_19(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_196_to_197),
    .west_valid_i          (valid_196_to_197),
    .west_ready_o          (ready_197_to_196),
    .west_data_o           (data_197_to_196),
    .west_valid_o          (valid_197_to_196),
    .west_ready_i          (ready_196_to_197),
    .east_data_i           (data_198_to_197),
    .east_valid_i          (valid_198_to_197),
    .east_ready_o          (ready_197_to_198),
    .east_data_o           (data_197_to_198),
    .east_valid_o          (valid_197_to_198),
    .east_ready_i          (ready_198_to_197),
    .vert0_data_i          (data_187_to_197_v0),
    .vert0_valid_i         (valid_187_to_197_v0),
    .vert0_ready_o         (ready_197_to_187_v0),
    .vert0_data_o          (data_197_to_207_v0),
    .vert0_valid_o         (valid_197_to_207_v0),
    .vert0_ready_i         (ready_207_to_197_v0),
    .vert1_data_i          (data_187_to_197_v1),
    .vert1_valid_i         (valid_187_to_197_v1),
    .vert1_ready_o         (ready_197_to_187_v1),
    .vert1_data_o          (data_197_to_207_v1),
    .vert1_valid_o         (valid_197_to_207_v1),
    .vert1_ready_i         (ready_207_to_197_v1),
    .local_data_i          (data_i[7][19]),
    .local_valid_i         (valid_i[7][19]),
    .local_ready_o         (ready_o[7][19]),
    .local_data_o          (data_o[7][19]),
    .local_valid_o         (valid_o[7][19]),
    .local_ready_i         (ready_i[7][19]),
    .credit_upd            (credit_upd)
);

/*Router 7,20*/    
cast_router #(
    .isUBM_list            (isUBM_list_7_20),
    .isFC_list             (isFC_list_7_20),
    .FCdn_list             (FCdn_list_7_20),
    .FCpl_list             (FCpl_list_7_20),
    .rt_file_list          (cast_rt_file_list_7_20)
)router_7_20(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_206_to_207),
    .west_valid_i          (valid_206_to_207),
    .west_ready_o          (ready_207_to_206),
    .west_data_o           (data_207_to_206),
    .west_valid_o          (valid_207_to_206),
    .west_ready_i          (ready_206_to_207),
    .east_data_i           (data_208_to_207),
    .east_valid_i          (valid_208_to_207),
    .east_ready_o          (ready_207_to_208),
    .east_data_o           (data_207_to_208),
    .east_valid_o          (valid_207_to_208),
    .east_ready_i          (ready_208_to_207),
    .vert0_data_i          (data_197_to_207_v0),
    .vert0_valid_i         (valid_197_to_207_v0),
    .vert0_ready_o         (ready_207_to_197_v0),
    .vert0_data_o          (data_207_to_217_v0),
    .vert0_valid_o         (valid_207_to_217_v0),
    .vert0_ready_i         (ready_217_to_207_v0),
    .vert1_data_i          (data_197_to_207_v1),
    .vert1_valid_i         (valid_197_to_207_v1),
    .vert1_ready_o         (ready_207_to_197_v1),
    .vert1_data_o          (data_207_to_217_v1),
    .vert1_valid_o         (valid_207_to_217_v1),
    .vert1_ready_i         (ready_217_to_207_v1),
    .local_data_i          (data_i[7][20]),
    .local_valid_i         (valid_i[7][20]),
    .local_ready_o         (ready_o[7][20]),
    .local_data_o          (data_o[7][20]),
    .local_valid_o         (valid_o[7][20]),
    .local_ready_i         (ready_i[7][20]),
    .credit_upd            (credit_upd)
);

/*Router 7,21*/    
cast_router #(
    .isUBM_list            (isUBM_list_7_21),
    .isFC_list             (isFC_list_7_21),
    .FCdn_list             (FCdn_list_7_21),
    .FCpl_list             (FCpl_list_7_21),
    .rt_file_list          (cast_rt_file_list_7_21)
)router_7_21(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_216_to_217),
    .west_valid_i          (valid_216_to_217),
    .west_ready_o          (ready_217_to_216),
    .west_data_o           (data_217_to_216),
    .west_valid_o          (valid_217_to_216),
    .west_ready_i          (ready_216_to_217),
    .east_data_i           (data_218_to_217),
    .east_valid_i          (valid_218_to_217),
    .east_ready_o          (ready_217_to_218),
    .east_data_o           (data_217_to_218),
    .east_valid_o          (valid_217_to_218),
    .east_ready_i          (ready_218_to_217),
    .vert0_data_i          (data_207_to_217_v0),
    .vert0_valid_i         (valid_207_to_217_v0),
    .vert0_ready_o         (ready_217_to_207_v0),
    .vert0_data_o          (data_217_to_227_v0),
    .vert0_valid_o         (valid_217_to_227_v0),
    .vert0_ready_i         (ready_227_to_217_v0),
    .vert1_data_i          (data_207_to_217_v1),
    .vert1_valid_i         (valid_207_to_217_v1),
    .vert1_ready_o         (ready_217_to_207_v1),
    .vert1_data_o          (data_217_to_227_v1),
    .vert1_valid_o         (valid_217_to_227_v1),
    .vert1_ready_i         (ready_227_to_217_v1),
    .local_data_i          (data_i[7][21]),
    .local_valid_i         (valid_i[7][21]),
    .local_ready_o         (ready_o[7][21]),
    .local_data_o          (data_o[7][21]),
    .local_valid_o         (valid_o[7][21]),
    .local_ready_i         (ready_i[7][21]),
    .credit_upd            (credit_upd)
);

/*Router 7,22*/    
cast_router #(
    .isUBM_list            (isUBM_list_7_22),
    .isFC_list             (isFC_list_7_22),
    .FCdn_list             (FCdn_list_7_22),
    .FCpl_list             (FCpl_list_7_22),
    .rt_file_list          (cast_rt_file_list_7_22)
)router_7_22(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_226_to_227),
    .west_valid_i          (valid_226_to_227),
    .west_ready_o          (ready_227_to_226),
    .west_data_o           (data_o_flee0),
    .west_valid_o          (valid_o_flee0),
    .west_ready_i          (ready_i_flee0),
    .east_data_i           (data_228_to_227),
    .east_valid_i          (valid_228_to_227),
    .east_ready_o          (ready_227_to_228),
    .east_data_o           (data_227_to_228),
    .east_valid_o          (valid_227_to_228),
    .east_ready_i          (ready_228_to_227),
    .vert0_data_i          (data_217_to_227_v0),
    .vert0_valid_i         (valid_217_to_227_v0),
    .vert0_ready_o         (ready_227_to_217_v0),
    .vert0_data_o          (data_227_to_237_v0),
    .vert0_valid_o         (valid_227_to_237_v0),
    .vert0_ready_i         (ready_237_to_227_v0),
    .vert1_data_i          (data_217_to_227_v1),
    .vert1_valid_i         (valid_217_to_227_v1),
    .vert1_ready_o         (ready_227_to_217_v1),
    .vert1_data_o          (data_227_to_237_v1),
    .vert1_valid_o         (valid_227_to_237_v1),
    .vert1_ready_i         (ready_237_to_227_v1),
    .local_data_i          (data_i[7][22]),
    .local_valid_i         (valid_i[7][22]),
    .local_ready_o         (ready_o[7][22]),
    .local_data_o          (data_o[7][22]),
    .local_valid_o         (valid_o[7][22]),
    .local_ready_i         (ready_i[7][22]),
    .credit_upd            (credit_upd)
);

/*Router 7,23*/    
cast_router #(
    .isUBM_list            (isUBM_list_7_23),
    .isFC_list             (isFC_list_7_23),
    .FCdn_list             (FCdn_list_7_23),
    .FCpl_list             (FCpl_list_7_23),
    .rt_file_list          (cast_rt_file_list_7_23)
)router_7_23(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_236_to_237),
    .west_valid_i          (valid_236_to_237),
    .west_ready_o          (ready_237_to_236),
    .west_data_o           (data_237_to_236),
    .west_valid_o          (valid_237_to_236),
    .west_ready_i          (ready_236_to_237),
    .east_data_i           (data_238_to_237),
    .east_valid_i          (valid_238_to_237),
    .east_ready_o          (ready_237_to_238),
    .east_data_o           (data_237_to_238),
    .east_valid_o          (valid_237_to_238),
    .east_ready_i          (ready_238_to_237),
    .vert0_data_i          (data_227_to_237_v0),
    .vert0_valid_i         (valid_227_to_237_v0),
    .vert0_ready_o         (ready_237_to_227_v0),
    .vert0_data_o          (data_237_to_247_v0),
    .vert0_valid_o         (valid_237_to_247_v0),
    .vert0_ready_i         (ready_247_to_237_v0),
    .vert1_data_i          (data_227_to_237_v1),
    .vert1_valid_i         (valid_227_to_237_v1),
    .vert1_ready_o         (ready_237_to_227_v1),
    .vert1_data_o          (data_237_to_247_v1),
    .vert1_valid_o         (valid_237_to_247_v1),
    .vert1_ready_i         (ready_247_to_237_v1),
    .local_data_i          (data_i[7][23]),
    .local_valid_i         (valid_i[7][23]),
    .local_ready_o         (ready_o[7][23]),
    .local_data_o          (data_o[7][23]),
    .local_valid_o         (valid_o[7][23]),
    .local_ready_i         (ready_i[7][23]),
    .credit_upd            (credit_upd)
);

/*Router 7,24*/    
cast_router #(
    .isUBM_list            (isUBM_list_7_24),
    .isFC_list             (isFC_list_7_24),
    .FCdn_list             (FCdn_list_7_24),
    .FCpl_list             (FCpl_list_7_24),
    .rt_file_list          (cast_rt_file_list_7_24)
)router_7_24(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_246_to_247),
    .west_valid_i          (valid_246_to_247),
    .west_ready_o          (ready_247_to_246),
    .west_data_o           (data_247_to_246),
    .west_valid_o          (valid_247_to_246),
    .west_ready_i          (ready_246_to_247),
    .east_data_i           (data_248_to_247),
    .east_valid_i          (valid_248_to_247),
    .east_ready_o          (ready_247_to_248),
    .east_data_o           (data_247_to_248),
    .east_valid_o          (valid_247_to_248),
    .east_ready_i          (ready_248_to_247),
    .vert0_data_i          (data_237_to_247_v0),
    .vert0_valid_i         (valid_237_to_247_v0),
    .vert0_ready_o         (ready_247_to_237_v0),
    .vert0_data_o          (),
    .vert0_valid_o         (),
    .vert0_ready_i         (1'b0),
    .vert1_data_i          (data_237_to_247_v1),
    .vert1_valid_i         (valid_237_to_247_v1),
    .vert1_ready_o         (ready_247_to_237_v1),
    .vert1_data_o          (),
    .vert1_valid_o         (),
    .vert1_ready_i         (1'b0),
    .local_data_i          (data_i[7][24]),
    .local_valid_i         (valid_i[7][24]),
    .local_ready_o         (ready_o[7][24]),
    .local_data_o          (data_o[7][24]),
    .local_valid_o         (valid_o[7][24]),
    .local_ready_i         (ready_i[7][24]),
    .credit_upd            (credit_upd)
);

/*Router 8,0*/    
cast_router #(
    .isUBM_list            (isUBM_list_8_0),
    .isFC_list             (isFC_list_8_0),
    .FCdn_list             (FCdn_list_8_0),
    .FCpl_list             (FCpl_list_8_0),
    .rt_file_list          (cast_rt_file_list_8_0)
)router_8_0(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_7_to_8),
    .west_valid_i          (valid_7_to_8),
    .west_ready_o          (ready_8_to_7),
    .west_data_o           (data_8_to_7),
    .west_valid_o          (valid_8_to_7),
    .west_ready_i          (ready_7_to_8),
    .east_data_i           (data_9_to_8),
    .east_valid_i          (valid_9_to_8),
    .east_ready_o          (ready_8_to_9),
    .east_data_o           (data_8_to_9),
    .east_valid_o          (valid_8_to_9),
    .east_ready_i          (ready_9_to_8),
    .vert0_data_i          (34'b0),
    .vert0_valid_i         (1'b0),
    .vert0_ready_o         (),
    .vert0_data_o          (data_8_to_18_v0),
    .vert0_valid_o         (valid_8_to_18_v0),
    .vert0_ready_i         (ready_18_to_8_v0),
    .vert1_data_i          (34'b0),
    .vert1_valid_i         (1'b0),
    .vert1_ready_o         (),
    .vert1_data_o          (data_8_to_18_v1),
    .vert1_valid_o         (valid_8_to_18_v1),
    .vert1_ready_i         (ready_18_to_8_v1),
    .local_data_i          (data_i[8][0]),
    .local_valid_i         (valid_i[8][0]),
    .local_ready_o         (ready_o[8][0]),
    .local_data_o          (data_o[8][0]),
    .local_valid_o         (valid_o[8][0]),
    .local_ready_i         (ready_i[8][0]),
    .credit_upd            (credit_upd)
);

/*Router 8,1*/    
cast_router #(
    .isUBM_list            (isUBM_list_8_1),
    .isFC_list             (isFC_list_8_1),
    .FCdn_list             (FCdn_list_8_1),
    .FCpl_list             (FCpl_list_8_1),
    .rt_file_list          (cast_rt_file_list_8_1)
)router_8_1(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_17_to_18),
    .west_valid_i          (valid_17_to_18),
    .west_ready_o          (ready_18_to_17),
    .west_data_o           (data_18_to_17),
    .west_valid_o          (valid_18_to_17),
    .west_ready_i          (ready_17_to_18),
    .east_data_i           (data_19_to_18),
    .east_valid_i          (valid_19_to_18),
    .east_ready_o          (ready_18_to_19),
    .east_data_o           (data_18_to_19),
    .east_valid_o          (valid_18_to_19),
    .east_ready_i          (ready_19_to_18),
    .vert0_data_i          (data_8_to_18_v0),
    .vert0_valid_i         (valid_8_to_18_v0),
    .vert0_ready_o         (ready_18_to_8_v0),
    .vert0_data_o          (data_18_to_28_v0),
    .vert0_valid_o         (valid_18_to_28_v0),
    .vert0_ready_i         (ready_28_to_18_v0),
    .vert1_data_i          (data_8_to_18_v1),
    .vert1_valid_i         (valid_8_to_18_v1),
    .vert1_ready_o         (ready_18_to_8_v1),
    .vert1_data_o          (data_18_to_28_v1),
    .vert1_valid_o         (valid_18_to_28_v1),
    .vert1_ready_i         (ready_28_to_18_v1),
    .local_data_i          (data_i[8][1]),
    .local_valid_i         (valid_i[8][1]),
    .local_ready_o         (ready_o[8][1]),
    .local_data_o          (data_o[8][1]),
    .local_valid_o         (valid_o[8][1]),
    .local_ready_i         (ready_i[8][1]),
    .credit_upd            (credit_upd)
);

/*Router 8,2*/    
cast_router #(
    .isUBM_list            (isUBM_list_8_2),
    .isFC_list             (isFC_list_8_2),
    .FCdn_list             (FCdn_list_8_2),
    .FCpl_list             (FCpl_list_8_2),
    .rt_file_list          (cast_rt_file_list_8_2)
)router_8_2(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_27_to_28),
    .west_valid_i          (valid_27_to_28),
    .west_ready_o          (ready_28_to_27),
    .west_data_o           (data_28_to_27),
    .west_valid_o          (valid_28_to_27),
    .west_ready_i          (ready_27_to_28),
    .east_data_i           (data_29_to_28),
    .east_valid_i          (valid_29_to_28),
    .east_ready_o          (ready_28_to_29),
    .east_data_o           (data_28_to_29),
    .east_valid_o          (valid_28_to_29),
    .east_ready_i          (ready_29_to_28),
    .vert0_data_i          (data_18_to_28_v0),
    .vert0_valid_i         (valid_18_to_28_v0),
    .vert0_ready_o         (ready_28_to_18_v0),
    .vert0_data_o          (data_28_to_38_v0),
    .vert0_valid_o         (valid_28_to_38_v0),
    .vert0_ready_i         (ready_38_to_28_v0),
    .vert1_data_i          (data_18_to_28_v1),
    .vert1_valid_i         (valid_18_to_28_v1),
    .vert1_ready_o         (ready_28_to_18_v1),
    .vert1_data_o          (data_28_to_38_v1),
    .vert1_valid_o         (valid_28_to_38_v1),
    .vert1_ready_i         (ready_38_to_28_v1),
    .local_data_i          (data_i[8][2]),
    .local_valid_i         (valid_i[8][2]),
    .local_ready_o         (ready_o[8][2]),
    .local_data_o          (data_o[8][2]),
    .local_valid_o         (valid_o[8][2]),
    .local_ready_i         (ready_i[8][2]),
    .credit_upd            (credit_upd)
);

/*Router 8,3*/    
cast_router #(
    .isUBM_list            (isUBM_list_8_3),
    .isFC_list             (isFC_list_8_3),
    .FCdn_list             (FCdn_list_8_3),
    .FCpl_list             (FCpl_list_8_3),
    .rt_file_list          (cast_rt_file_list_8_3)
)router_8_3(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_37_to_38),
    .west_valid_i          (valid_37_to_38),
    .west_ready_o          (ready_38_to_37),
    .west_data_o           (data_38_to_37),
    .west_valid_o          (valid_38_to_37),
    .west_ready_i          (ready_37_to_38),
    .east_data_i           (data_39_to_38),
    .east_valid_i          (valid_39_to_38),
    .east_ready_o          (ready_38_to_39),
    .east_data_o           (data_38_to_39),
    .east_valid_o          (valid_38_to_39),
    .east_ready_i          (ready_39_to_38),
    .vert0_data_i          (data_28_to_38_v0),
    .vert0_valid_i         (valid_28_to_38_v0),
    .vert0_ready_o         (ready_38_to_28_v0),
    .vert0_data_o          (data_38_to_48_v0),
    .vert0_valid_o         (valid_38_to_48_v0),
    .vert0_ready_i         (ready_48_to_38_v0),
    .vert1_data_i          (data_28_to_38_v1),
    .vert1_valid_i         (valid_28_to_38_v1),
    .vert1_ready_o         (ready_38_to_28_v1),
    .vert1_data_o          (data_38_to_48_v1),
    .vert1_valid_o         (valid_38_to_48_v1),
    .vert1_ready_i         (ready_48_to_38_v1),
    .local_data_i          (data_i[8][3]),
    .local_valid_i         (valid_i[8][3]),
    .local_ready_o         (ready_o[8][3]),
    .local_data_o          (data_o[8][3]),
    .local_valid_o         (valid_o[8][3]),
    .local_ready_i         (ready_i[8][3]),
    .credit_upd            (credit_upd)
);

/*Router 8,4*/    
cast_router #(
    .isUBM_list            (isUBM_list_8_4),
    .isFC_list             (isFC_list_8_4),
    .FCdn_list             (FCdn_list_8_4),
    .FCpl_list             (FCpl_list_8_4),
    .rt_file_list          (cast_rt_file_list_8_4)
)router_8_4(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_47_to_48),
    .west_valid_i          (valid_47_to_48),
    .west_ready_o          (ready_48_to_47),
    .west_data_o           (data_48_to_47),
    .west_valid_o          (valid_48_to_47),
    .west_ready_i          (ready_47_to_48),
    .east_data_i           (data_49_to_48),
    .east_valid_i          (valid_49_to_48),
    .east_ready_o          (ready_48_to_49),
    .east_data_o           (data_48_to_49),
    .east_valid_o          (valid_48_to_49),
    .east_ready_i          (ready_49_to_48),
    .vert0_data_i          (data_38_to_48_v0),
    .vert0_valid_i         (valid_38_to_48_v0),
    .vert0_ready_o         (ready_48_to_38_v0),
    .vert0_data_o          (data_48_to_58_v0),
    .vert0_valid_o         (valid_48_to_58_v0),
    .vert0_ready_i         (ready_58_to_48_v0),
    .vert1_data_i          (data_38_to_48_v1),
    .vert1_valid_i         (valid_38_to_48_v1),
    .vert1_ready_o         (ready_48_to_38_v1),
    .vert1_data_o          (data_48_to_58_v1),
    .vert1_valid_o         (valid_48_to_58_v1),
    .vert1_ready_i         (ready_58_to_48_v1),
    .local_data_i          (data_i[8][4]),
    .local_valid_i         (valid_i[8][4]),
    .local_ready_o         (ready_o[8][4]),
    .local_data_o          (data_o[8][4]),
    .local_valid_o         (valid_o[8][4]),
    .local_ready_i         (ready_i[8][4]),
    .credit_upd            (credit_upd)
);

/*Router 8,5*/    
cast_router #(
    .isUBM_list            (isUBM_list_8_5),
    .isFC_list             (isFC_list_8_5),
    .FCdn_list             (FCdn_list_8_5),
    .FCpl_list             (FCpl_list_8_5),
    .rt_file_list          (cast_rt_file_list_8_5)
)router_8_5(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_57_to_58),
    .west_valid_i          (valid_57_to_58),
    .west_ready_o          (ready_58_to_57),
    .west_data_o           (data_58_to_57),
    .west_valid_o          (valid_58_to_57),
    .west_ready_i          (ready_57_to_58),
    .east_data_i           (data_59_to_58),
    .east_valid_i          (valid_59_to_58),
    .east_ready_o          (ready_58_to_59),
    .east_data_o           (data_58_to_59),
    .east_valid_o          (valid_58_to_59),
    .east_ready_i          (ready_59_to_58),
    .vert0_data_i          (data_48_to_58_v0),
    .vert0_valid_i         (valid_48_to_58_v0),
    .vert0_ready_o         (ready_58_to_48_v0),
    .vert0_data_o          (data_58_to_68_v0),
    .vert0_valid_o         (valid_58_to_68_v0),
    .vert0_ready_i         (ready_68_to_58_v0),
    .vert1_data_i          (data_48_to_58_v1),
    .vert1_valid_i         (valid_48_to_58_v1),
    .vert1_ready_o         (ready_58_to_48_v1),
    .vert1_data_o          (data_58_to_68_v1),
    .vert1_valid_o         (valid_58_to_68_v1),
    .vert1_ready_i         (ready_68_to_58_v1),
    .local_data_i          (data_i[8][5]),
    .local_valid_i         (valid_i[8][5]),
    .local_ready_o         (ready_o[8][5]),
    .local_data_o          (data_o[8][5]),
    .local_valid_o         (valid_o[8][5]),
    .local_ready_i         (ready_i[8][5]),
    .credit_upd            (credit_upd)
);

/*Router 8,6*/    
cast_router #(
    .isUBM_list            (isUBM_list_8_6),
    .isFC_list             (isFC_list_8_6),
    .FCdn_list             (FCdn_list_8_6),
    .FCpl_list             (FCpl_list_8_6),
    .rt_file_list          (cast_rt_file_list_8_6)
)router_8_6(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_67_to_68),
    .west_valid_i          (valid_67_to_68),
    .west_ready_o          (ready_68_to_67),
    .west_data_o           (data_68_to_67),
    .west_valid_o          (valid_68_to_67),
    .west_ready_i          (ready_67_to_68),
    .east_data_i           (data_69_to_68),
    .east_valid_i          (valid_69_to_68),
    .east_ready_o          (ready_68_to_69),
    .east_data_o           (data_68_to_69),
    .east_valid_o          (valid_68_to_69),
    .east_ready_i          (ready_69_to_68),
    .vert0_data_i          (data_58_to_68_v0),
    .vert0_valid_i         (valid_58_to_68_v0),
    .vert0_ready_o         (ready_68_to_58_v0),
    .vert0_data_o          (data_68_to_78_v0),
    .vert0_valid_o         (valid_68_to_78_v0),
    .vert0_ready_i         (ready_78_to_68_v0),
    .vert1_data_i          (data_58_to_68_v1),
    .vert1_valid_i         (valid_58_to_68_v1),
    .vert1_ready_o         (ready_68_to_58_v1),
    .vert1_data_o          (data_68_to_78_v1),
    .vert1_valid_o         (valid_68_to_78_v1),
    .vert1_ready_i         (ready_78_to_68_v1),
    .local_data_i          (data_i[8][6]),
    .local_valid_i         (valid_i[8][6]),
    .local_ready_o         (ready_o[8][6]),
    .local_data_o          (data_o[8][6]),
    .local_valid_o         (valid_o[8][6]),
    .local_ready_i         (ready_i[8][6]),
    .credit_upd            (credit_upd)
);

/*Router 8,7*/    
cast_router #(
    .isUBM_list            (isUBM_list_8_7),
    .isFC_list             (isFC_list_8_7),
    .FCdn_list             (FCdn_list_8_7),
    .FCpl_list             (FCpl_list_8_7),
    .rt_file_list          (cast_rt_file_list_8_7)
)router_8_7(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_77_to_78),
    .west_valid_i          (valid_77_to_78),
    .west_ready_o          (ready_78_to_77),
    .west_data_o           (data_78_to_77),
    .west_valid_o          (valid_78_to_77),
    .west_ready_i          (ready_77_to_78),
    .east_data_i           (data_79_to_78),
    .east_valid_i          (valid_79_to_78),
    .east_ready_o          (ready_78_to_79),
    .east_data_o           (data_78_to_79),
    .east_valid_o          (valid_78_to_79),
    .east_ready_i          (ready_79_to_78),
    .vert0_data_i          (data_68_to_78_v0),
    .vert0_valid_i         (valid_68_to_78_v0),
    .vert0_ready_o         (ready_78_to_68_v0),
    .vert0_data_o          (data_78_to_88_v0),
    .vert0_valid_o         (valid_78_to_88_v0),
    .vert0_ready_i         (ready_88_to_78_v0),
    .vert1_data_i          (data_68_to_78_v1),
    .vert1_valid_i         (valid_68_to_78_v1),
    .vert1_ready_o         (ready_78_to_68_v1),
    .vert1_data_o          (data_78_to_88_v1),
    .vert1_valid_o         (valid_78_to_88_v1),
    .vert1_ready_i         (ready_88_to_78_v1),
    .local_data_i          (data_i[8][7]),
    .local_valid_i         (valid_i[8][7]),
    .local_ready_o         (ready_o[8][7]),
    .local_data_o          (data_o[8][7]),
    .local_valid_o         (valid_o[8][7]),
    .local_ready_i         (ready_i[8][7]),
    .credit_upd            (credit_upd)
);

/*Router 8,8*/    
cast_router #(
    .isUBM_list            (isUBM_list_8_8),
    .isFC_list             (isFC_list_8_8),
    .FCdn_list             (FCdn_list_8_8),
    .FCpl_list             (FCpl_list_8_8),
    .rt_file_list          (cast_rt_file_list_8_8)
)router_8_8(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_87_to_88),
    .west_valid_i          (valid_87_to_88),
    .west_ready_o          (ready_88_to_87),
    .west_data_o           (data_88_to_87),
    .west_valid_o          (valid_88_to_87),
    .west_ready_i          (ready_87_to_88),
    .east_data_i           (data_89_to_88),
    .east_valid_i          (valid_89_to_88),
    .east_ready_o          (ready_88_to_89),
    .east_data_o           (data_88_to_89),
    .east_valid_o          (valid_88_to_89),
    .east_ready_i          (ready_89_to_88),
    .vert0_data_i          (data_78_to_88_v0),
    .vert0_valid_i         (valid_78_to_88_v0),
    .vert0_ready_o         (ready_88_to_78_v0),
    .vert0_data_o          (data_88_to_98_v0),
    .vert0_valid_o         (valid_88_to_98_v0),
    .vert0_ready_i         (ready_98_to_88_v0),
    .vert1_data_i          (data_78_to_88_v1),
    .vert1_valid_i         (valid_78_to_88_v1),
    .vert1_ready_o         (ready_88_to_78_v1),
    .vert1_data_o          (data_88_to_98_v1),
    .vert1_valid_o         (valid_88_to_98_v1),
    .vert1_ready_i         (ready_98_to_88_v1),
    .local_data_i          (data_i[8][8]),
    .local_valid_i         (valid_i[8][8]),
    .local_ready_o         (ready_o[8][8]),
    .local_data_o          (data_o[8][8]),
    .local_valid_o         (valid_o[8][8]),
    .local_ready_i         (ready_i[8][8]),
    .credit_upd            (credit_upd)
);

/*Router 8,9*/    
cast_router #(
    .isUBM_list            (isUBM_list_8_9),
    .isFC_list             (isFC_list_8_9),
    .FCdn_list             (FCdn_list_8_9),
    .FCpl_list             (FCpl_list_8_9),
    .rt_file_list          (cast_rt_file_list_8_9)
)router_8_9(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_97_to_98),
    .west_valid_i          (valid_97_to_98),
    .west_ready_o          (ready_98_to_97),
    .west_data_o           (data_98_to_97),
    .west_valid_o          (valid_98_to_97),
    .west_ready_i          (ready_97_to_98),
    .east_data_i           (data_99_to_98),
    .east_valid_i          (valid_99_to_98),
    .east_ready_o          (ready_98_to_99),
    .east_data_o           (data_98_to_99),
    .east_valid_o          (valid_98_to_99),
    .east_ready_i          (ready_99_to_98),
    .vert0_data_i          (data_88_to_98_v0),
    .vert0_valid_i         (valid_88_to_98_v0),
    .vert0_ready_o         (ready_98_to_88_v0),
    .vert0_data_o          (data_98_to_108_v0),
    .vert0_valid_o         (valid_98_to_108_v0),
    .vert0_ready_i         (ready_108_to_98_v0),
    .vert1_data_i          (data_88_to_98_v1),
    .vert1_valid_i         (valid_88_to_98_v1),
    .vert1_ready_o         (ready_98_to_88_v1),
    .vert1_data_o          (data_98_to_108_v1),
    .vert1_valid_o         (valid_98_to_108_v1),
    .vert1_ready_i         (ready_108_to_98_v1),
    .local_data_i          (data_i[8][9]),
    .local_valid_i         (valid_i[8][9]),
    .local_ready_o         (ready_o[8][9]),
    .local_data_o          (data_o[8][9]),
    .local_valid_o         (valid_o[8][9]),
    .local_ready_i         (ready_i[8][9]),
    .credit_upd            (credit_upd)
);

/*Router 8,10*/    
cast_router #(
    .isUBM_list            (isUBM_list_8_10),
    .isFC_list             (isFC_list_8_10),
    .FCdn_list             (FCdn_list_8_10),
    .FCpl_list             (FCpl_list_8_10),
    .rt_file_list          (cast_rt_file_list_8_10)
)router_8_10(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_107_to_108),
    .west_valid_i          (valid_107_to_108),
    .west_ready_o          (ready_108_to_107),
    .west_data_o           (data_108_to_107),
    .west_valid_o          (valid_108_to_107),
    .west_ready_i          (ready_107_to_108),
    .east_data_i           (data_109_to_108),
    .east_valid_i          (valid_109_to_108),
    .east_ready_o          (ready_108_to_109),
    .east_data_o           (data_108_to_109),
    .east_valid_o          (valid_108_to_109),
    .east_ready_i          (ready_109_to_108),
    .vert0_data_i          (data_98_to_108_v0),
    .vert0_valid_i         (valid_98_to_108_v0),
    .vert0_ready_o         (ready_108_to_98_v0),
    .vert0_data_o          (data_108_to_118_v0),
    .vert0_valid_o         (valid_108_to_118_v0),
    .vert0_ready_i         (ready_118_to_108_v0),
    .vert1_data_i          (data_98_to_108_v1),
    .vert1_valid_i         (valid_98_to_108_v1),
    .vert1_ready_o         (ready_108_to_98_v1),
    .vert1_data_o          (data_108_to_118_v1),
    .vert1_valid_o         (valid_108_to_118_v1),
    .vert1_ready_i         (ready_118_to_108_v1),
    .local_data_i          (data_i[8][10]),
    .local_valid_i         (valid_i[8][10]),
    .local_ready_o         (ready_o[8][10]),
    .local_data_o          (data_o[8][10]),
    .local_valid_o         (valid_o[8][10]),
    .local_ready_i         (ready_i[8][10]),
    .credit_upd            (credit_upd)
);

/*Router 8,11*/    
cast_router #(
    .isUBM_list            (isUBM_list_8_11),
    .isFC_list             (isFC_list_8_11),
    .FCdn_list             (FCdn_list_8_11),
    .FCpl_list             (FCpl_list_8_11),
    .rt_file_list          (cast_rt_file_list_8_11)
)router_8_11(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_117_to_118),
    .west_valid_i          (valid_117_to_118),
    .west_ready_o          (ready_118_to_117),
    .west_data_o           (data_118_to_117),
    .west_valid_o          (valid_118_to_117),
    .west_ready_i          (ready_117_to_118),
    .east_data_i           (data_119_to_118),
    .east_valid_i          (valid_119_to_118),
    .east_ready_o          (ready_118_to_119),
    .east_data_o           (data_118_to_119),
    .east_valid_o          (valid_118_to_119),
    .east_ready_i          (ready_119_to_118),
    .vert0_data_i          (data_108_to_118_v0),
    .vert0_valid_i         (valid_108_to_118_v0),
    .vert0_ready_o         (ready_118_to_108_v0),
    .vert0_data_o          (data_118_to_128_v0),
    .vert0_valid_o         (valid_118_to_128_v0),
    .vert0_ready_i         (ready_128_to_118_v0),
    .vert1_data_i          (data_108_to_118_v1),
    .vert1_valid_i         (valid_108_to_118_v1),
    .vert1_ready_o         (ready_118_to_108_v1),
    .vert1_data_o          (data_118_to_128_v1),
    .vert1_valid_o         (valid_118_to_128_v1),
    .vert1_ready_i         (ready_128_to_118_v1),
    .local_data_i          (data_i[8][11]),
    .local_valid_i         (valid_i[8][11]),
    .local_ready_o         (ready_o[8][11]),
    .local_data_o          (data_o[8][11]),
    .local_valid_o         (valid_o[8][11]),
    .local_ready_i         (ready_i[8][11]),
    .credit_upd            (credit_upd)
);

/*Router 8,12*/    
cast_router #(
    .isUBM_list            (isUBM_list_8_12),
    .isFC_list             (isFC_list_8_12),
    .FCdn_list             (FCdn_list_8_12),
    .FCpl_list             (FCpl_list_8_12),
    .rt_file_list          (cast_rt_file_list_8_12)
)router_8_12(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_127_to_128),
    .west_valid_i          (valid_127_to_128),
    .west_ready_o          (ready_128_to_127),
    .west_data_o           (data_128_to_127),
    .west_valid_o          (valid_128_to_127),
    .west_ready_i          (ready_127_to_128),
    .east_data_i           (data_129_to_128),
    .east_valid_i          (valid_129_to_128),
    .east_ready_o          (ready_128_to_129),
    .east_data_o           (data_128_to_129),
    .east_valid_o          (valid_128_to_129),
    .east_ready_i          (ready_129_to_128),
    .vert0_data_i          (data_118_to_128_v0),
    .vert0_valid_i         (valid_118_to_128_v0),
    .vert0_ready_o         (ready_128_to_118_v0),
    .vert0_data_o          (data_128_to_138_v0),
    .vert0_valid_o         (valid_128_to_138_v0),
    .vert0_ready_i         (ready_138_to_128_v0),
    .vert1_data_i          (data_118_to_128_v1),
    .vert1_valid_i         (valid_118_to_128_v1),
    .vert1_ready_o         (ready_128_to_118_v1),
    .vert1_data_o          (data_128_to_138_v1),
    .vert1_valid_o         (valid_128_to_138_v1),
    .vert1_ready_i         (ready_138_to_128_v1),
    .local_data_i          (data_i[8][12]),
    .local_valid_i         (valid_i[8][12]),
    .local_ready_o         (ready_o[8][12]),
    .local_data_o          (data_o[8][12]),
    .local_valid_o         (valid_o[8][12]),
    .local_ready_i         (ready_i[8][12]),
    .credit_upd            (credit_upd)
);

/*Router 8,13*/    
cast_router #(
    .isUBM_list            (isUBM_list_8_13),
    .isFC_list             (isFC_list_8_13),
    .FCdn_list             (FCdn_list_8_13),
    .FCpl_list             (FCpl_list_8_13),
    .rt_file_list          (cast_rt_file_list_8_13)
)router_8_13(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_137_to_138),
    .west_valid_i          (valid_137_to_138),
    .west_ready_o          (ready_138_to_137),
    .west_data_o           (data_138_to_137),
    .west_valid_o          (valid_138_to_137),
    .west_ready_i          (ready_137_to_138),
    .east_data_i           (data_139_to_138),
    .east_valid_i          (valid_139_to_138),
    .east_ready_o          (ready_138_to_139),
    .east_data_o           (data_138_to_139),
    .east_valid_o          (valid_138_to_139),
    .east_ready_i          (ready_139_to_138),
    .vert0_data_i          (data_128_to_138_v0),
    .vert0_valid_i         (valid_128_to_138_v0),
    .vert0_ready_o         (ready_138_to_128_v0),
    .vert0_data_o          (data_138_to_148_v0),
    .vert0_valid_o         (valid_138_to_148_v0),
    .vert0_ready_i         (ready_148_to_138_v0),
    .vert1_data_i          (data_128_to_138_v1),
    .vert1_valid_i         (valid_128_to_138_v1),
    .vert1_ready_o         (ready_138_to_128_v1),
    .vert1_data_o          (data_138_to_148_v1),
    .vert1_valid_o         (valid_138_to_148_v1),
    .vert1_ready_i         (ready_148_to_138_v1),
    .local_data_i          (data_i[8][13]),
    .local_valid_i         (valid_i[8][13]),
    .local_ready_o         (ready_o[8][13]),
    .local_data_o          (data_o[8][13]),
    .local_valid_o         (valid_o[8][13]),
    .local_ready_i         (ready_i[8][13]),
    .credit_upd            (credit_upd)
);

/*Router 8,14*/    
cast_router #(
    .isUBM_list            (isUBM_list_8_14),
    .isFC_list             (isFC_list_8_14),
    .FCdn_list             (FCdn_list_8_14),
    .FCpl_list             (FCpl_list_8_14),
    .rt_file_list          (cast_rt_file_list_8_14)
)router_8_14(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_147_to_148),
    .west_valid_i          (valid_147_to_148),
    .west_ready_o          (ready_148_to_147),
    .west_data_o           (data_148_to_147),
    .west_valid_o          (valid_148_to_147),
    .west_ready_i          (ready_147_to_148),
    .east_data_i           (data_149_to_148),
    .east_valid_i          (valid_149_to_148),
    .east_ready_o          (ready_148_to_149),
    .east_data_o           (data_148_to_149),
    .east_valid_o          (valid_148_to_149),
    .east_ready_i          (ready_149_to_148),
    .vert0_data_i          (data_138_to_148_v0),
    .vert0_valid_i         (valid_138_to_148_v0),
    .vert0_ready_o         (ready_148_to_138_v0),
    .vert0_data_o          (data_148_to_158_v0),
    .vert0_valid_o         (valid_148_to_158_v0),
    .vert0_ready_i         (ready_158_to_148_v0),
    .vert1_data_i          (data_138_to_148_v1),
    .vert1_valid_i         (valid_138_to_148_v1),
    .vert1_ready_o         (ready_148_to_138_v1),
    .vert1_data_o          (data_148_to_158_v1),
    .vert1_valid_o         (valid_148_to_158_v1),
    .vert1_ready_i         (ready_158_to_148_v1),
    .local_data_i          (data_i[8][14]),
    .local_valid_i         (valid_i[8][14]),
    .local_ready_o         (ready_o[8][14]),
    .local_data_o          (data_o[8][14]),
    .local_valid_o         (valid_o[8][14]),
    .local_ready_i         (ready_i[8][14]),
    .credit_upd            (credit_upd)
);

/*Router 8,15*/    
cast_router #(
    .isUBM_list            (isUBM_list_8_15),
    .isFC_list             (isFC_list_8_15),
    .FCdn_list             (FCdn_list_8_15),
    .FCpl_list             (FCpl_list_8_15),
    .rt_file_list          (cast_rt_file_list_8_15)
)router_8_15(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_157_to_158),
    .west_valid_i          (valid_157_to_158),
    .west_ready_o          (ready_158_to_157),
    .west_data_o           (data_158_to_157),
    .west_valid_o          (valid_158_to_157),
    .west_ready_i          (ready_157_to_158),
    .east_data_i           (data_159_to_158),
    .east_valid_i          (valid_159_to_158),
    .east_ready_o          (ready_158_to_159),
    .east_data_o           (data_158_to_159),
    .east_valid_o          (valid_158_to_159),
    .east_ready_i          (ready_159_to_158),
    .vert0_data_i          (data_148_to_158_v0),
    .vert0_valid_i         (valid_148_to_158_v0),
    .vert0_ready_o         (ready_158_to_148_v0),
    .vert0_data_o          (data_158_to_168_v0),
    .vert0_valid_o         (valid_158_to_168_v0),
    .vert0_ready_i         (ready_168_to_158_v0),
    .vert1_data_i          (data_148_to_158_v1),
    .vert1_valid_i         (valid_148_to_158_v1),
    .vert1_ready_o         (ready_158_to_148_v1),
    .vert1_data_o          (data_158_to_168_v1),
    .vert1_valid_o         (valid_158_to_168_v1),
    .vert1_ready_i         (ready_168_to_158_v1),
    .local_data_i          (data_i[8][15]),
    .local_valid_i         (valid_i[8][15]),
    .local_ready_o         (ready_o[8][15]),
    .local_data_o          (data_o[8][15]),
    .local_valid_o         (valid_o[8][15]),
    .local_ready_i         (ready_i[8][15]),
    .credit_upd            (credit_upd)
);

/*Router 8,16*/    
cast_router #(
    .isUBM_list            (isUBM_list_8_16),
    .isFC_list             (isFC_list_8_16),
    .FCdn_list             (FCdn_list_8_16),
    .FCpl_list             (FCpl_list_8_16),
    .rt_file_list          (cast_rt_file_list_8_16)
)router_8_16(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_167_to_168),
    .west_valid_i          (valid_167_to_168),
    .west_ready_o          (ready_168_to_167),
    .west_data_o           (data_168_to_167),
    .west_valid_o          (valid_168_to_167),
    .west_ready_i          (ready_167_to_168),
    .east_data_i           (data_169_to_168),
    .east_valid_i          (valid_169_to_168),
    .east_ready_o          (ready_168_to_169),
    .east_data_o           (data_168_to_169),
    .east_valid_o          (valid_168_to_169),
    .east_ready_i          (ready_169_to_168),
    .vert0_data_i          (data_158_to_168_v0),
    .vert0_valid_i         (valid_158_to_168_v0),
    .vert0_ready_o         (ready_168_to_158_v0),
    .vert0_data_o          (data_168_to_178_v0),
    .vert0_valid_o         (valid_168_to_178_v0),
    .vert0_ready_i         (ready_178_to_168_v0),
    .vert1_data_i          (data_158_to_168_v1),
    .vert1_valid_i         (valid_158_to_168_v1),
    .vert1_ready_o         (ready_168_to_158_v1),
    .vert1_data_o          (data_168_to_178_v1),
    .vert1_valid_o         (valid_168_to_178_v1),
    .vert1_ready_i         (ready_178_to_168_v1),
    .local_data_i          (data_i[8][16]),
    .local_valid_i         (valid_i[8][16]),
    .local_ready_o         (ready_o[8][16]),
    .local_data_o          (data_o[8][16]),
    .local_valid_o         (valid_o[8][16]),
    .local_ready_i         (ready_i[8][16]),
    .credit_upd            (credit_upd)
);

/*Router 8,17*/    
cast_router #(
    .isUBM_list            (isUBM_list_8_17),
    .isFC_list             (isFC_list_8_17),
    .FCdn_list             (FCdn_list_8_17),
    .FCpl_list             (FCpl_list_8_17),
    .rt_file_list          (cast_rt_file_list_8_17)
)router_8_17(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_177_to_178),
    .west_valid_i          (valid_177_to_178),
    .west_ready_o          (ready_178_to_177),
    .west_data_o           (data_178_to_177),
    .west_valid_o          (valid_178_to_177),
    .west_ready_i          (ready_177_to_178),
    .east_data_i           (data_179_to_178),
    .east_valid_i          (valid_179_to_178),
    .east_ready_o          (ready_178_to_179),
    .east_data_o           (data_178_to_179),
    .east_valid_o          (valid_178_to_179),
    .east_ready_i          (ready_179_to_178),
    .vert0_data_i          (data_168_to_178_v0),
    .vert0_valid_i         (valid_168_to_178_v0),
    .vert0_ready_o         (ready_178_to_168_v0),
    .vert0_data_o          (data_178_to_188_v0),
    .vert0_valid_o         (valid_178_to_188_v0),
    .vert0_ready_i         (ready_188_to_178_v0),
    .vert1_data_i          (data_168_to_178_v1),
    .vert1_valid_i         (valid_168_to_178_v1),
    .vert1_ready_o         (ready_178_to_168_v1),
    .vert1_data_o          (data_178_to_188_v1),
    .vert1_valid_o         (valid_178_to_188_v1),
    .vert1_ready_i         (ready_188_to_178_v1),
    .local_data_i          (data_i[8][17]),
    .local_valid_i         (valid_i[8][17]),
    .local_ready_o         (ready_o[8][17]),
    .local_data_o          (data_o[8][17]),
    .local_valid_o         (valid_o[8][17]),
    .local_ready_i         (ready_i[8][17]),
    .credit_upd            (credit_upd)
);

/*Router 8,18*/    
cast_router #(
    .isUBM_list            (isUBM_list_8_18),
    .isFC_list             (isFC_list_8_18),
    .FCdn_list             (FCdn_list_8_18),
    .FCpl_list             (FCpl_list_8_18),
    .rt_file_list          (cast_rt_file_list_8_18)
)router_8_18(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_187_to_188),
    .west_valid_i          (valid_187_to_188),
    .west_ready_o          (ready_188_to_187),
    .west_data_o           (data_188_to_187),
    .west_valid_o          (valid_188_to_187),
    .west_ready_i          (ready_187_to_188),
    .east_data_i           (data_189_to_188),
    .east_valid_i          (valid_189_to_188),
    .east_ready_o          (ready_188_to_189),
    .east_data_o           (data_188_to_189),
    .east_valid_o          (valid_188_to_189),
    .east_ready_i          (ready_189_to_188),
    .vert0_data_i          (data_178_to_188_v0),
    .vert0_valid_i         (valid_178_to_188_v0),
    .vert0_ready_o         (ready_188_to_178_v0),
    .vert0_data_o          (data_188_to_198_v0),
    .vert0_valid_o         (valid_188_to_198_v0),
    .vert0_ready_i         (ready_198_to_188_v0),
    .vert1_data_i          (data_178_to_188_v1),
    .vert1_valid_i         (valid_178_to_188_v1),
    .vert1_ready_o         (ready_188_to_178_v1),
    .vert1_data_o          (data_188_to_198_v1),
    .vert1_valid_o         (valid_188_to_198_v1),
    .vert1_ready_i         (ready_198_to_188_v1),
    .local_data_i          (data_i[8][18]),
    .local_valid_i         (valid_i[8][18]),
    .local_ready_o         (ready_o[8][18]),
    .local_data_o          (data_o[8][18]),
    .local_valid_o         (valid_o[8][18]),
    .local_ready_i         (ready_i[8][18]),
    .credit_upd            (credit_upd)
);

/*Router 8,19*/    
cast_router #(
    .isUBM_list            (isUBM_list_8_19),
    .isFC_list             (isFC_list_8_19),
    .FCdn_list             (FCdn_list_8_19),
    .FCpl_list             (FCpl_list_8_19),
    .rt_file_list          (cast_rt_file_list_8_19)
)router_8_19(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_197_to_198),
    .west_valid_i          (valid_197_to_198),
    .west_ready_o          (ready_198_to_197),
    .west_data_o           (data_198_to_197),
    .west_valid_o          (valid_198_to_197),
    .west_ready_i          (ready_197_to_198),
    .east_data_i           (data_199_to_198),
    .east_valid_i          (valid_199_to_198),
    .east_ready_o          (ready_198_to_199),
    .east_data_o           (data_198_to_199),
    .east_valid_o          (valid_198_to_199),
    .east_ready_i          (ready_199_to_198),
    .vert0_data_i          (data_188_to_198_v0),
    .vert0_valid_i         (valid_188_to_198_v0),
    .vert0_ready_o         (ready_198_to_188_v0),
    .vert0_data_o          (data_198_to_208_v0),
    .vert0_valid_o         (valid_198_to_208_v0),
    .vert0_ready_i         (ready_208_to_198_v0),
    .vert1_data_i          (data_188_to_198_v1),
    .vert1_valid_i         (valid_188_to_198_v1),
    .vert1_ready_o         (ready_198_to_188_v1),
    .vert1_data_o          (data_198_to_208_v1),
    .vert1_valid_o         (valid_198_to_208_v1),
    .vert1_ready_i         (ready_208_to_198_v1),
    .local_data_i          (data_i[8][19]),
    .local_valid_i         (valid_i[8][19]),
    .local_ready_o         (ready_o[8][19]),
    .local_data_o          (data_o[8][19]),
    .local_valid_o         (valid_o[8][19]),
    .local_ready_i         (ready_i[8][19]),
    .credit_upd            (credit_upd)
);

/*Router 8,20*/    
cast_router #(
    .isUBM_list            (isUBM_list_8_20),
    .isFC_list             (isFC_list_8_20),
    .FCdn_list             (FCdn_list_8_20),
    .FCpl_list             (FCpl_list_8_20),
    .rt_file_list          (cast_rt_file_list_8_20)
)router_8_20(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_207_to_208),
    .west_valid_i          (valid_207_to_208),
    .west_ready_o          (ready_208_to_207),
    .west_data_o           (data_208_to_207),
    .west_valid_o          (valid_208_to_207),
    .west_ready_i          (ready_207_to_208),
    .east_data_i           (data_209_to_208),
    .east_valid_i          (valid_209_to_208),
    .east_ready_o          (ready_208_to_209),
    .east_data_o           (data_208_to_209),
    .east_valid_o          (valid_208_to_209),
    .east_ready_i          (ready_209_to_208),
    .vert0_data_i          (data_198_to_208_v0),
    .vert0_valid_i         (valid_198_to_208_v0),
    .vert0_ready_o         (ready_208_to_198_v0),
    .vert0_data_o          (data_208_to_218_v0),
    .vert0_valid_o         (valid_208_to_218_v0),
    .vert0_ready_i         (ready_218_to_208_v0),
    .vert1_data_i          (data_198_to_208_v1),
    .vert1_valid_i         (valid_198_to_208_v1),
    .vert1_ready_o         (ready_208_to_198_v1),
    .vert1_data_o          (data_208_to_218_v1),
    .vert1_valid_o         (valid_208_to_218_v1),
    .vert1_ready_i         (ready_218_to_208_v1),
    .local_data_i          (data_i[8][20]),
    .local_valid_i         (valid_i[8][20]),
    .local_ready_o         (ready_o[8][20]),
    .local_data_o          (data_o[8][20]),
    .local_valid_o         (valid_o[8][20]),
    .local_ready_i         (ready_i[8][20]),
    .credit_upd            (credit_upd)
);

/*Router 8,21*/    
cast_router #(
    .isUBM_list            (isUBM_list_8_21),
    .isFC_list             (isFC_list_8_21),
    .FCdn_list             (FCdn_list_8_21),
    .FCpl_list             (FCpl_list_8_21),
    .rt_file_list          (cast_rt_file_list_8_21)
)router_8_21(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_217_to_218),
    .west_valid_i          (valid_217_to_218),
    .west_ready_o          (ready_218_to_217),
    .west_data_o           (data_218_to_217),
    .west_valid_o          (valid_218_to_217),
    .west_ready_i          (ready_217_to_218),
    .east_data_i           (data_219_to_218),
    .east_valid_i          (valid_219_to_218),
    .east_ready_o          (ready_218_to_219),
    .east_data_o           (data_218_to_219),
    .east_valid_o          (valid_218_to_219),
    .east_ready_i          (ready_219_to_218),
    .vert0_data_i          (data_208_to_218_v0),
    .vert0_valid_i         (valid_208_to_218_v0),
    .vert0_ready_o         (ready_218_to_208_v0),
    .vert0_data_o          (data_218_to_228_v0),
    .vert0_valid_o         (valid_218_to_228_v0),
    .vert0_ready_i         (ready_228_to_218_v0),
    .vert1_data_i          (data_208_to_218_v1),
    .vert1_valid_i         (valid_208_to_218_v1),
    .vert1_ready_o         (ready_218_to_208_v1),
    .vert1_data_o          (data_218_to_228_v1),
    .vert1_valid_o         (valid_218_to_228_v1),
    .vert1_ready_i         (ready_228_to_218_v1),
    .local_data_i          (data_i[8][21]),
    .local_valid_i         (valid_i[8][21]),
    .local_ready_o         (ready_o[8][21]),
    .local_data_o          (data_o[8][21]),
    .local_valid_o         (valid_o[8][21]),
    .local_ready_i         (ready_i[8][21]),
    .credit_upd            (credit_upd)
);

/*Router 8,22*/    
cast_router #(
    .isUBM_list            (isUBM_list_8_22),
    .isFC_list             (isFC_list_8_22),
    .FCdn_list             (FCdn_list_8_22),
    .FCpl_list             (FCpl_list_8_22),
    .rt_file_list          (cast_rt_file_list_8_22)
)router_8_22(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_227_to_228),
    .west_valid_i          (valid_227_to_228),
    .west_ready_o          (ready_228_to_227),
    .west_data_o           (data_228_to_227),
    .west_valid_o          (valid_228_to_227),
    .west_ready_i          (ready_227_to_228),
    .east_data_i           (data_229_to_228),
    .east_valid_i          (valid_229_to_228),
    .east_ready_o          (ready_228_to_229),
    .east_data_o           (data_228_to_229),
    .east_valid_o          (valid_228_to_229),
    .east_ready_i          (ready_229_to_228),
    .vert0_data_i          (data_218_to_228_v0),
    .vert0_valid_i         (valid_218_to_228_v0),
    .vert0_ready_o         (ready_228_to_218_v0),
    .vert0_data_o          (data_228_to_238_v0),
    .vert0_valid_o         (valid_228_to_238_v0),
    .vert0_ready_i         (ready_238_to_228_v0),
    .vert1_data_i          (data_218_to_228_v1),
    .vert1_valid_i         (valid_218_to_228_v1),
    .vert1_ready_o         (ready_228_to_218_v1),
    .vert1_data_o          (data_228_to_238_v1),
    .vert1_valid_o         (valid_228_to_238_v1),
    .vert1_ready_i         (ready_238_to_228_v1),
    .local_data_i          (data_i[8][22]),
    .local_valid_i         (valid_i[8][22]),
    .local_ready_o         (ready_o[8][22]),
    .local_data_o          (data_o[8][22]),
    .local_valid_o         (valid_o[8][22]),
    .local_ready_i         (ready_i[8][22]),
    .credit_upd            (credit_upd)
);

/*Router 8,23*/    
cast_router #(
    .isUBM_list            (isUBM_list_8_23),
    .isFC_list             (isFC_list_8_23),
    .FCdn_list             (FCdn_list_8_23),
    .FCpl_list             (FCpl_list_8_23),
    .rt_file_list          (cast_rt_file_list_8_23)
)router_8_23(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_237_to_238),
    .west_valid_i          (valid_237_to_238),
    .west_ready_o          (ready_238_to_237),
    .west_data_o           (data_o_flee2),
    .west_valid_o          (valid_o_flee2),
    .west_ready_i          (ready_i_flee2),
    .east_data_i           (data_239_to_238),
    .east_valid_i          (valid_239_to_238),
    .east_ready_o          (ready_238_to_239),
    .east_data_o           (data_238_to_239),
    .east_valid_o          (valid_238_to_239),
    .east_ready_i          (ready_239_to_238),
    .vert0_data_i          (data_228_to_238_v0),
    .vert0_valid_i         (valid_228_to_238_v0),
    .vert0_ready_o         (ready_238_to_228_v0),
    .vert0_data_o          (data_238_to_248_v0),
    .vert0_valid_o         (valid_238_to_248_v0),
    .vert0_ready_i         (ready_248_to_238_v0),
    .vert1_data_i          (data_228_to_238_v1),
    .vert1_valid_i         (valid_228_to_238_v1),
    .vert1_ready_o         (ready_238_to_228_v1),
    .vert1_data_o          (data_238_to_248_v1),
    .vert1_valid_o         (valid_238_to_248_v1),
    .vert1_ready_i         (ready_248_to_238_v1),
    .local_data_i          (data_i[8][23]),
    .local_valid_i         (valid_i[8][23]),
    .local_ready_o         (ready_o[8][23]),
    .local_data_o          (data_o[8][23]),
    .local_valid_o         (valid_o[8][23]),
    .local_ready_i         (ready_i[8][23]),
    .credit_upd            (credit_upd)
);

/*Router 8,24*/    
cast_router #(
    .isUBM_list            (isUBM_list_8_24),
    .isFC_list             (isFC_list_8_24),
    .FCdn_list             (FCdn_list_8_24),
    .FCpl_list             (FCpl_list_8_24),
    .rt_file_list          (cast_rt_file_list_8_24)
)router_8_24(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_247_to_248),
    .west_valid_i          (valid_247_to_248),
    .west_ready_o          (ready_248_to_247),
    .west_data_o           (data_248_to_247),
    .west_valid_o          (valid_248_to_247),
    .west_ready_i          (ready_247_to_248),
    .east_data_i           (data_249_to_248),
    .east_valid_i          (valid_249_to_248),
    .east_ready_o          (ready_248_to_249),
    .east_data_o           (data_248_to_249),
    .east_valid_o          (valid_248_to_249),
    .east_ready_i          (ready_249_to_248),
    .vert0_data_i          (data_238_to_248_v0),
    .vert0_valid_i         (valid_238_to_248_v0),
    .vert0_ready_o         (ready_248_to_238_v0),
    .vert0_data_o          (),
    .vert0_valid_o         (),
    .vert0_ready_i         (1'b0),
    .vert1_data_i          (data_238_to_248_v1),
    .vert1_valid_i         (valid_238_to_248_v1),
    .vert1_ready_o         (ready_248_to_238_v1),
    .vert1_data_o          (),
    .vert1_valid_o         (),
    .vert1_ready_i         (1'b0),
    .local_data_i          (data_i[8][24]),
    .local_valid_i         (valid_i[8][24]),
    .local_ready_o         (ready_o[8][24]),
    .local_data_o          (data_o[8][24]),
    .local_valid_o         (valid_o[8][24]),
    .local_ready_i         (ready_i[8][24]),
    .credit_upd            (credit_upd)
);

/*Router 9,0*/    
cast_router #(
    .isUBM_list            (isUBM_list_9_0),
    .isFC_list             (isFC_list_9_0),
    .FCdn_list             (FCdn_list_9_0),
    .FCpl_list             (FCpl_list_9_0),
    .rt_file_list          (cast_rt_file_list_9_0)
)router_9_0(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_8_to_9),
    .west_valid_i          (valid_8_to_9),
    .west_ready_o          (ready_9_to_8),
    .west_data_o           (data_9_to_8),
    .west_valid_o          (valid_9_to_8),
    .west_ready_i          (ready_8_to_9),
    .east_data_i           (34'b0),
    .east_valid_i          (1'b0),
    .east_ready_o          (),
    .east_data_o           (),
    .east_valid_o          (),
    .east_ready_i          (1'b0),
    .vert0_data_i          (34'b0),
    .vert0_valid_i         (1'b0),
    .vert0_ready_o         (),
    .vert0_data_o          (data_9_to_19_v0),
    .vert0_valid_o         (valid_9_to_19_v0),
    .vert0_ready_i         (ready_19_to_9_v0),
    .vert1_data_i          (34'b0),
    .vert1_valid_i         (1'b0),
    .vert1_ready_o         (),
    .vert1_data_o          (data_9_to_19_v1),
    .vert1_valid_o         (valid_9_to_19_v1),
    .vert1_ready_i         (ready_19_to_9_v1),
    .local_data_i          (data_i[9][0]),
    .local_valid_i         (valid_i[9][0]),
    .local_ready_o         (ready_o[9][0]),
    .local_data_o          (data_o[9][0]),
    .local_valid_o         (valid_o[9][0]),
    .local_ready_i         (ready_i[9][0]),
    .credit_upd            (credit_upd)
);

/*Router 9,1*/    
cast_router #(
    .isUBM_list            (isUBM_list_9_1),
    .isFC_list             (isFC_list_9_1),
    .FCdn_list             (FCdn_list_9_1),
    .FCpl_list             (FCpl_list_9_1),
    .rt_file_list          (cast_rt_file_list_9_1)
)router_9_1(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_18_to_19),
    .west_valid_i          (valid_18_to_19),
    .west_ready_o          (ready_19_to_18),
    .west_data_o           (data_19_to_18),
    .west_valid_o          (valid_19_to_18),
    .west_ready_i          (ready_18_to_19),
    .east_data_i           (34'b0),
    .east_valid_i          (1'b0),
    .east_ready_o          (),
    .east_data_o           (),
    .east_valid_o          (),
    .east_ready_i          (1'b0),
    .vert0_data_i          (data_9_to_19_v0),
    .vert0_valid_i         (valid_9_to_19_v0),
    .vert0_ready_o         (ready_19_to_9_v0),
    .vert0_data_o          (data_19_to_29_v0),
    .vert0_valid_o         (valid_19_to_29_v0),
    .vert0_ready_i         (ready_29_to_19_v0),
    .vert1_data_i          (data_9_to_19_v1),
    .vert1_valid_i         (valid_9_to_19_v1),
    .vert1_ready_o         (ready_19_to_9_v1),
    .vert1_data_o          (data_19_to_29_v1),
    .vert1_valid_o         (valid_19_to_29_v1),
    .vert1_ready_i         (ready_29_to_19_v1),
    .local_data_i          (data_i[9][1]),
    .local_valid_i         (valid_i[9][1]),
    .local_ready_o         (ready_o[9][1]),
    .local_data_o          (data_o[9][1]),
    .local_valid_o         (valid_o[9][1]),
    .local_ready_i         (ready_i[9][1]),
    .credit_upd            (credit_upd)
);

/*Router 9,2*/    
cast_router #(
    .isUBM_list            (isUBM_list_9_2),
    .isFC_list             (isFC_list_9_2),
    .FCdn_list             (FCdn_list_9_2),
    .FCpl_list             (FCpl_list_9_2),
    .rt_file_list          (cast_rt_file_list_9_2)
)router_9_2(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_28_to_29),
    .west_valid_i          (valid_28_to_29),
    .west_ready_o          (ready_29_to_28),
    .west_data_o           (data_29_to_28),
    .west_valid_o          (valid_29_to_28),
    .west_ready_i          (ready_28_to_29),
    .east_data_i           (34'b0),
    .east_valid_i          (1'b0),
    .east_ready_o          (),
    .east_data_o           (),
    .east_valid_o          (),
    .east_ready_i          (1'b0),
    .vert0_data_i          (data_19_to_29_v0),
    .vert0_valid_i         (valid_19_to_29_v0),
    .vert0_ready_o         (ready_29_to_19_v0),
    .vert0_data_o          (data_29_to_39_v0),
    .vert0_valid_o         (valid_29_to_39_v0),
    .vert0_ready_i         (ready_39_to_29_v0),
    .vert1_data_i          (data_19_to_29_v1),
    .vert1_valid_i         (valid_19_to_29_v1),
    .vert1_ready_o         (ready_29_to_19_v1),
    .vert1_data_o          (data_29_to_39_v1),
    .vert1_valid_o         (valid_29_to_39_v1),
    .vert1_ready_i         (ready_39_to_29_v1),
    .local_data_i          (data_i[9][2]),
    .local_valid_i         (valid_i[9][2]),
    .local_ready_o         (ready_o[9][2]),
    .local_data_o          (data_o[9][2]),
    .local_valid_o         (valid_o[9][2]),
    .local_ready_i         (ready_i[9][2]),
    .credit_upd            (credit_upd)
);

/*Router 9,3*/    
cast_router #(
    .isUBM_list            (isUBM_list_9_3),
    .isFC_list             (isFC_list_9_3),
    .FCdn_list             (FCdn_list_9_3),
    .FCpl_list             (FCpl_list_9_3),
    .rt_file_list          (cast_rt_file_list_9_3)
)router_9_3(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_38_to_39),
    .west_valid_i          (valid_38_to_39),
    .west_ready_o          (ready_39_to_38),
    .west_data_o           (data_39_to_38),
    .west_valid_o          (valid_39_to_38),
    .west_ready_i          (ready_38_to_39),
    .east_data_i           (34'b0),
    .east_valid_i          (1'b0),
    .east_ready_o          (),
    .east_data_o           (),
    .east_valid_o          (),
    .east_ready_i          (1'b0),
    .vert0_data_i          (data_29_to_39_v0),
    .vert0_valid_i         (valid_29_to_39_v0),
    .vert0_ready_o         (ready_39_to_29_v0),
    .vert0_data_o          (data_39_to_49_v0),
    .vert0_valid_o         (valid_39_to_49_v0),
    .vert0_ready_i         (ready_49_to_39_v0),
    .vert1_data_i          (data_29_to_39_v1),
    .vert1_valid_i         (valid_29_to_39_v1),
    .vert1_ready_o         (ready_39_to_29_v1),
    .vert1_data_o          (data_39_to_49_v1),
    .vert1_valid_o         (valid_39_to_49_v1),
    .vert1_ready_i         (ready_49_to_39_v1),
    .local_data_i          (data_i[9][3]),
    .local_valid_i         (valid_i[9][3]),
    .local_ready_o         (ready_o[9][3]),
    .local_data_o          (data_o[9][3]),
    .local_valid_o         (valid_o[9][3]),
    .local_ready_i         (ready_i[9][3]),
    .credit_upd            (credit_upd)
);

/*Router 9,4*/    
cast_router #(
    .isUBM_list            (isUBM_list_9_4),
    .isFC_list             (isFC_list_9_4),
    .FCdn_list             (FCdn_list_9_4),
    .FCpl_list             (FCpl_list_9_4),
    .rt_file_list          (cast_rt_file_list_9_4)
)router_9_4(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_48_to_49),
    .west_valid_i          (valid_48_to_49),
    .west_ready_o          (ready_49_to_48),
    .west_data_o           (data_49_to_48),
    .west_valid_o          (valid_49_to_48),
    .west_ready_i          (ready_48_to_49),
    .east_data_i           (34'b0),
    .east_valid_i          (1'b0),
    .east_ready_o          (),
    .east_data_o           (),
    .east_valid_o          (),
    .east_ready_i          (1'b0),
    .vert0_data_i          (data_39_to_49_v0),
    .vert0_valid_i         (valid_39_to_49_v0),
    .vert0_ready_o         (ready_49_to_39_v0),
    .vert0_data_o          (data_49_to_59_v0),
    .vert0_valid_o         (valid_49_to_59_v0),
    .vert0_ready_i         (ready_59_to_49_v0),
    .vert1_data_i          (data_39_to_49_v1),
    .vert1_valid_i         (valid_39_to_49_v1),
    .vert1_ready_o         (ready_49_to_39_v1),
    .vert1_data_o          (data_49_to_59_v1),
    .vert1_valid_o         (valid_49_to_59_v1),
    .vert1_ready_i         (ready_59_to_49_v1),
    .local_data_i          (data_i[9][4]),
    .local_valid_i         (valid_i[9][4]),
    .local_ready_o         (ready_o[9][4]),
    .local_data_o          (data_o[9][4]),
    .local_valid_o         (valid_o[9][4]),
    .local_ready_i         (ready_i[9][4]),
    .credit_upd            (credit_upd)
);

/*Router 9,5*/    
cast_router #(
    .isUBM_list            (isUBM_list_9_5),
    .isFC_list             (isFC_list_9_5),
    .FCdn_list             (FCdn_list_9_5),
    .FCpl_list             (FCpl_list_9_5),
    .rt_file_list          (cast_rt_file_list_9_5)
)router_9_5(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_58_to_59),
    .west_valid_i          (valid_58_to_59),
    .west_ready_o          (ready_59_to_58),
    .west_data_o           (data_59_to_58),
    .west_valid_o          (valid_59_to_58),
    .west_ready_i          (ready_58_to_59),
    .east_data_i           (34'b0),
    .east_valid_i          (1'b0),
    .east_ready_o          (),
    .east_data_o           (),
    .east_valid_o          (),
    .east_ready_i          (1'b0),
    .vert0_data_i          (data_49_to_59_v0),
    .vert0_valid_i         (valid_49_to_59_v0),
    .vert0_ready_o         (ready_59_to_49_v0),
    .vert0_data_o          (data_59_to_69_v0),
    .vert0_valid_o         (valid_59_to_69_v0),
    .vert0_ready_i         (ready_69_to_59_v0),
    .vert1_data_i          (data_49_to_59_v1),
    .vert1_valid_i         (valid_49_to_59_v1),
    .vert1_ready_o         (ready_59_to_49_v1),
    .vert1_data_o          (data_59_to_69_v1),
    .vert1_valid_o         (valid_59_to_69_v1),
    .vert1_ready_i         (ready_69_to_59_v1),
    .local_data_i          (data_i[9][5]),
    .local_valid_i         (valid_i[9][5]),
    .local_ready_o         (ready_o[9][5]),
    .local_data_o          (data_o[9][5]),
    .local_valid_o         (valid_o[9][5]),
    .local_ready_i         (ready_i[9][5]),
    .credit_upd            (credit_upd)
);

/*Router 9,6*/    
cast_router #(
    .isUBM_list            (isUBM_list_9_6),
    .isFC_list             (isFC_list_9_6),
    .FCdn_list             (FCdn_list_9_6),
    .FCpl_list             (FCpl_list_9_6),
    .rt_file_list          (cast_rt_file_list_9_6)
)router_9_6(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_68_to_69),
    .west_valid_i          (valid_68_to_69),
    .west_ready_o          (ready_69_to_68),
    .west_data_o           (data_69_to_68),
    .west_valid_o          (valid_69_to_68),
    .west_ready_i          (ready_68_to_69),
    .east_data_i           (34'b0),
    .east_valid_i          (1'b0),
    .east_ready_o          (),
    .east_data_o           (),
    .east_valid_o          (),
    .east_ready_i          (1'b0),
    .vert0_data_i          (data_59_to_69_v0),
    .vert0_valid_i         (valid_59_to_69_v0),
    .vert0_ready_o         (ready_69_to_59_v0),
    .vert0_data_o          (data_69_to_79_v0),
    .vert0_valid_o         (valid_69_to_79_v0),
    .vert0_ready_i         (ready_79_to_69_v0),
    .vert1_data_i          (data_59_to_69_v1),
    .vert1_valid_i         (valid_59_to_69_v1),
    .vert1_ready_o         (ready_69_to_59_v1),
    .vert1_data_o          (data_69_to_79_v1),
    .vert1_valid_o         (valid_69_to_79_v1),
    .vert1_ready_i         (ready_79_to_69_v1),
    .local_data_i          (data_i[9][6]),
    .local_valid_i         (valid_i[9][6]),
    .local_ready_o         (ready_o[9][6]),
    .local_data_o          (data_o[9][6]),
    .local_valid_o         (valid_o[9][6]),
    .local_ready_i         (ready_i[9][6]),
    .credit_upd            (credit_upd)
);

/*Router 9,7*/    
cast_router #(
    .isUBM_list            (isUBM_list_9_7),
    .isFC_list             (isFC_list_9_7),
    .FCdn_list             (FCdn_list_9_7),
    .FCpl_list             (FCpl_list_9_7),
    .rt_file_list          (cast_rt_file_list_9_7)
)router_9_7(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_78_to_79),
    .west_valid_i          (valid_78_to_79),
    .west_ready_o          (ready_79_to_78),
    .west_data_o           (data_79_to_78),
    .west_valid_o          (valid_79_to_78),
    .west_ready_i          (ready_78_to_79),
    .east_data_i           (34'b0),
    .east_valid_i          (1'b0),
    .east_ready_o          (),
    .east_data_o           (),
    .east_valid_o          (),
    .east_ready_i          (1'b0),
    .vert0_data_i          (data_69_to_79_v0),
    .vert0_valid_i         (valid_69_to_79_v0),
    .vert0_ready_o         (ready_79_to_69_v0),
    .vert0_data_o          (data_79_to_89_v0),
    .vert0_valid_o         (valid_79_to_89_v0),
    .vert0_ready_i         (ready_89_to_79_v0),
    .vert1_data_i          (data_69_to_79_v1),
    .vert1_valid_i         (valid_69_to_79_v1),
    .vert1_ready_o         (ready_79_to_69_v1),
    .vert1_data_o          (data_79_to_89_v1),
    .vert1_valid_o         (valid_79_to_89_v1),
    .vert1_ready_i         (ready_89_to_79_v1),
    .local_data_i          (data_i[9][7]),
    .local_valid_i         (valid_i[9][7]),
    .local_ready_o         (ready_o[9][7]),
    .local_data_o          (data_o[9][7]),
    .local_valid_o         (valid_o[9][7]),
    .local_ready_i         (ready_i[9][7]),
    .credit_upd            (credit_upd)
);

/*Router 9,8*/    
cast_router #(
    .isUBM_list            (isUBM_list_9_8),
    .isFC_list             (isFC_list_9_8),
    .FCdn_list             (FCdn_list_9_8),
    .FCpl_list             (FCpl_list_9_8),
    .rt_file_list          (cast_rt_file_list_9_8)
)router_9_8(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_88_to_89),
    .west_valid_i          (valid_88_to_89),
    .west_ready_o          (ready_89_to_88),
    .west_data_o           (data_89_to_88),
    .west_valid_o          (valid_89_to_88),
    .west_ready_i          (ready_88_to_89),
    .east_data_i           (34'b0),
    .east_valid_i          (1'b0),
    .east_ready_o          (),
    .east_data_o           (),
    .east_valid_o          (),
    .east_ready_i          (1'b0),
    .vert0_data_i          (data_79_to_89_v0),
    .vert0_valid_i         (valid_79_to_89_v0),
    .vert0_ready_o         (ready_89_to_79_v0),
    .vert0_data_o          (data_89_to_99_v0),
    .vert0_valid_o         (valid_89_to_99_v0),
    .vert0_ready_i         (ready_99_to_89_v0),
    .vert1_data_i          (data_79_to_89_v1),
    .vert1_valid_i         (valid_79_to_89_v1),
    .vert1_ready_o         (ready_89_to_79_v1),
    .vert1_data_o          (data_89_to_99_v1),
    .vert1_valid_o         (valid_89_to_99_v1),
    .vert1_ready_i         (ready_99_to_89_v1),
    .local_data_i          (data_i[9][8]),
    .local_valid_i         (valid_i[9][8]),
    .local_ready_o         (ready_o[9][8]),
    .local_data_o          (data_o[9][8]),
    .local_valid_o         (valid_o[9][8]),
    .local_ready_i         (ready_i[9][8]),
    .credit_upd            (credit_upd)
);

/*Router 9,9*/    
cast_router #(
    .isUBM_list            (isUBM_list_9_9),
    .isFC_list             (isFC_list_9_9),
    .FCdn_list             (FCdn_list_9_9),
    .FCpl_list             (FCpl_list_9_9),
    .rt_file_list          (cast_rt_file_list_9_9)
)router_9_9(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_98_to_99),
    .west_valid_i          (valid_98_to_99),
    .west_ready_o          (ready_99_to_98),
    .west_data_o           (data_99_to_98),
    .west_valid_o          (valid_99_to_98),
    .west_ready_i          (ready_98_to_99),
    .east_data_i           (34'b0),
    .east_valid_i          (1'b0),
    .east_ready_o          (),
    .east_data_o           (),
    .east_valid_o          (),
    .east_ready_i          (1'b0),
    .vert0_data_i          (data_89_to_99_v0),
    .vert0_valid_i         (valid_89_to_99_v0),
    .vert0_ready_o         (ready_99_to_89_v0),
    .vert0_data_o          (data_99_to_109_v0),
    .vert0_valid_o         (valid_99_to_109_v0),
    .vert0_ready_i         (ready_109_to_99_v0),
    .vert1_data_i          (data_89_to_99_v1),
    .vert1_valid_i         (valid_89_to_99_v1),
    .vert1_ready_o         (ready_99_to_89_v1),
    .vert1_data_o          (data_99_to_109_v1),
    .vert1_valid_o         (valid_99_to_109_v1),
    .vert1_ready_i         (ready_109_to_99_v1),
    .local_data_i          (data_i[9][9]),
    .local_valid_i         (valid_i[9][9]),
    .local_ready_o         (ready_o[9][9]),
    .local_data_o          (data_o[9][9]),
    .local_valid_o         (valid_o[9][9]),
    .local_ready_i         (ready_i[9][9]),
    .credit_upd            (credit_upd)
);

/*Router 9,10*/    
cast_router #(
    .isUBM_list            (isUBM_list_9_10),
    .isFC_list             (isFC_list_9_10),
    .FCdn_list             (FCdn_list_9_10),
    .FCpl_list             (FCpl_list_9_10),
    .rt_file_list          (cast_rt_file_list_9_10)
)router_9_10(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_108_to_109),
    .west_valid_i          (valid_108_to_109),
    .west_ready_o          (ready_109_to_108),
    .west_data_o           (data_109_to_108),
    .west_valid_o          (valid_109_to_108),
    .west_ready_i          (ready_108_to_109),
    .east_data_i           (34'b0),
    .east_valid_i          (1'b0),
    .east_ready_o          (),
    .east_data_o           (),
    .east_valid_o          (),
    .east_ready_i          (1'b0),
    .vert0_data_i          (data_99_to_109_v0),
    .vert0_valid_i         (valid_99_to_109_v0),
    .vert0_ready_o         (ready_109_to_99_v0),
    .vert0_data_o          (data_109_to_119_v0),
    .vert0_valid_o         (valid_109_to_119_v0),
    .vert0_ready_i         (ready_119_to_109_v0),
    .vert1_data_i          (data_99_to_109_v1),
    .vert1_valid_i         (valid_99_to_109_v1),
    .vert1_ready_o         (ready_109_to_99_v1),
    .vert1_data_o          (data_109_to_119_v1),
    .vert1_valid_o         (valid_109_to_119_v1),
    .vert1_ready_i         (ready_119_to_109_v1),
    .local_data_i          (data_i[9][10]),
    .local_valid_i         (valid_i[9][10]),
    .local_ready_o         (ready_o[9][10]),
    .local_data_o          (data_o[9][10]),
    .local_valid_o         (valid_o[9][10]),
    .local_ready_i         (ready_i[9][10]),
    .credit_upd            (credit_upd)
);

/*Router 9,11*/    
cast_router #(
    .isUBM_list            (isUBM_list_9_11),
    .isFC_list             (isFC_list_9_11),
    .FCdn_list             (FCdn_list_9_11),
    .FCpl_list             (FCpl_list_9_11),
    .rt_file_list          (cast_rt_file_list_9_11)
)router_9_11(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_118_to_119),
    .west_valid_i          (valid_118_to_119),
    .west_ready_o          (ready_119_to_118),
    .west_data_o           (data_119_to_118),
    .west_valid_o          (valid_119_to_118),
    .west_ready_i          (ready_118_to_119),
    .east_data_i           (34'b0),
    .east_valid_i          (1'b0),
    .east_ready_o          (),
    .east_data_o           (),
    .east_valid_o          (),
    .east_ready_i          (1'b0),
    .vert0_data_i          (data_109_to_119_v0),
    .vert0_valid_i         (valid_109_to_119_v0),
    .vert0_ready_o         (ready_119_to_109_v0),
    .vert0_data_o          (data_119_to_129_v0),
    .vert0_valid_o         (valid_119_to_129_v0),
    .vert0_ready_i         (ready_129_to_119_v0),
    .vert1_data_i          (data_109_to_119_v1),
    .vert1_valid_i         (valid_109_to_119_v1),
    .vert1_ready_o         (ready_119_to_109_v1),
    .vert1_data_o          (data_119_to_129_v1),
    .vert1_valid_o         (valid_119_to_129_v1),
    .vert1_ready_i         (ready_129_to_119_v1),
    .local_data_i          (data_i[9][11]),
    .local_valid_i         (valid_i[9][11]),
    .local_ready_o         (ready_o[9][11]),
    .local_data_o          (data_o[9][11]),
    .local_valid_o         (valid_o[9][11]),
    .local_ready_i         (ready_i[9][11]),
    .credit_upd            (credit_upd)
);

/*Router 9,12*/    
cast_router #(
    .isUBM_list            (isUBM_list_9_12),
    .isFC_list             (isFC_list_9_12),
    .FCdn_list             (FCdn_list_9_12),
    .FCpl_list             (FCpl_list_9_12),
    .rt_file_list          (cast_rt_file_list_9_12)
)router_9_12(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_128_to_129),
    .west_valid_i          (valid_128_to_129),
    .west_ready_o          (ready_129_to_128),
    .west_data_o           (data_129_to_128),
    .west_valid_o          (valid_129_to_128),
    .west_ready_i          (ready_128_to_129),
    .east_data_i           (34'b0),
    .east_valid_i          (1'b0),
    .east_ready_o          (),
    .east_data_o           (),
    .east_valid_o          (),
    .east_ready_i          (1'b0),
    .vert0_data_i          (data_119_to_129_v0),
    .vert0_valid_i         (valid_119_to_129_v0),
    .vert0_ready_o         (ready_129_to_119_v0),
    .vert0_data_o          (data_129_to_139_v0),
    .vert0_valid_o         (valid_129_to_139_v0),
    .vert0_ready_i         (ready_139_to_129_v0),
    .vert1_data_i          (data_119_to_129_v1),
    .vert1_valid_i         (valid_119_to_129_v1),
    .vert1_ready_o         (ready_129_to_119_v1),
    .vert1_data_o          (data_129_to_139_v1),
    .vert1_valid_o         (valid_129_to_139_v1),
    .vert1_ready_i         (ready_139_to_129_v1),
    .local_data_i          (data_i[9][12]),
    .local_valid_i         (valid_i[9][12]),
    .local_ready_o         (ready_o[9][12]),
    .local_data_o          (data_o[9][12]),
    .local_valid_o         (valid_o[9][12]),
    .local_ready_i         (ready_i[9][12]),
    .credit_upd            (credit_upd)
);

/*Router 9,13*/    
cast_router #(
    .isUBM_list            (isUBM_list_9_13),
    .isFC_list             (isFC_list_9_13),
    .FCdn_list             (FCdn_list_9_13),
    .FCpl_list             (FCpl_list_9_13),
    .rt_file_list          (cast_rt_file_list_9_13)
)router_9_13(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_138_to_139),
    .west_valid_i          (valid_138_to_139),
    .west_ready_o          (ready_139_to_138),
    .west_data_o           (data_139_to_138),
    .west_valid_o          (valid_139_to_138),
    .west_ready_i          (ready_138_to_139),
    .east_data_i           (34'b0),
    .east_valid_i          (1'b0),
    .east_ready_o          (),
    .east_data_o           (),
    .east_valid_o          (),
    .east_ready_i          (1'b0),
    .vert0_data_i          (data_129_to_139_v0),
    .vert0_valid_i         (valid_129_to_139_v0),
    .vert0_ready_o         (ready_139_to_129_v0),
    .vert0_data_o          (data_139_to_149_v0),
    .vert0_valid_o         (valid_139_to_149_v0),
    .vert0_ready_i         (ready_149_to_139_v0),
    .vert1_data_i          (data_129_to_139_v1),
    .vert1_valid_i         (valid_129_to_139_v1),
    .vert1_ready_o         (ready_139_to_129_v1),
    .vert1_data_o          (data_139_to_149_v1),
    .vert1_valid_o         (valid_139_to_149_v1),
    .vert1_ready_i         (ready_149_to_139_v1),
    .local_data_i          (data_i[9][13]),
    .local_valid_i         (valid_i[9][13]),
    .local_ready_o         (ready_o[9][13]),
    .local_data_o          (data_o[9][13]),
    .local_valid_o         (valid_o[9][13]),
    .local_ready_i         (ready_i[9][13]),
    .credit_upd            (credit_upd)
);

/*Router 9,14*/    
cast_router #(
    .isUBM_list            (isUBM_list_9_14),
    .isFC_list             (isFC_list_9_14),
    .FCdn_list             (FCdn_list_9_14),
    .FCpl_list             (FCpl_list_9_14),
    .rt_file_list          (cast_rt_file_list_9_14)
)router_9_14(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_148_to_149),
    .west_valid_i          (valid_148_to_149),
    .west_ready_o          (ready_149_to_148),
    .west_data_o           (data_149_to_148),
    .west_valid_o          (valid_149_to_148),
    .west_ready_i          (ready_148_to_149),
    .east_data_i           (34'b0),
    .east_valid_i          (1'b0),
    .east_ready_o          (),
    .east_data_o           (),
    .east_valid_o          (),
    .east_ready_i          (1'b0),
    .vert0_data_i          (data_139_to_149_v0),
    .vert0_valid_i         (valid_139_to_149_v0),
    .vert0_ready_o         (ready_149_to_139_v0),
    .vert0_data_o          (data_149_to_159_v0),
    .vert0_valid_o         (valid_149_to_159_v0),
    .vert0_ready_i         (ready_159_to_149_v0),
    .vert1_data_i          (data_139_to_149_v1),
    .vert1_valid_i         (valid_139_to_149_v1),
    .vert1_ready_o         (ready_149_to_139_v1),
    .vert1_data_o          (data_149_to_159_v1),
    .vert1_valid_o         (valid_149_to_159_v1),
    .vert1_ready_i         (ready_159_to_149_v1),
    .local_data_i          (data_i[9][14]),
    .local_valid_i         (valid_i[9][14]),
    .local_ready_o         (ready_o[9][14]),
    .local_data_o          (data_o[9][14]),
    .local_valid_o         (valid_o[9][14]),
    .local_ready_i         (ready_i[9][14]),
    .credit_upd            (credit_upd)
);

/*Router 9,15*/    
cast_router #(
    .isUBM_list            (isUBM_list_9_15),
    .isFC_list             (isFC_list_9_15),
    .FCdn_list             (FCdn_list_9_15),
    .FCpl_list             (FCpl_list_9_15),
    .rt_file_list          (cast_rt_file_list_9_15)
)router_9_15(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_158_to_159),
    .west_valid_i          (valid_158_to_159),
    .west_ready_o          (ready_159_to_158),
    .west_data_o           (data_159_to_158),
    .west_valid_o          (valid_159_to_158),
    .west_ready_i          (ready_158_to_159),
    .east_data_i           (34'b0),
    .east_valid_i          (1'b0),
    .east_ready_o          (),
    .east_data_o           (),
    .east_valid_o          (),
    .east_ready_i          (1'b0),
    .vert0_data_i          (data_149_to_159_v0),
    .vert0_valid_i         (valid_149_to_159_v0),
    .vert0_ready_o         (ready_159_to_149_v0),
    .vert0_data_o          (data_159_to_169_v0),
    .vert0_valid_o         (valid_159_to_169_v0),
    .vert0_ready_i         (ready_169_to_159_v0),
    .vert1_data_i          (data_149_to_159_v1),
    .vert1_valid_i         (valid_149_to_159_v1),
    .vert1_ready_o         (ready_159_to_149_v1),
    .vert1_data_o          (data_159_to_169_v1),
    .vert1_valid_o         (valid_159_to_169_v1),
    .vert1_ready_i         (ready_169_to_159_v1),
    .local_data_i          (data_i[9][15]),
    .local_valid_i         (valid_i[9][15]),
    .local_ready_o         (ready_o[9][15]),
    .local_data_o          (data_o[9][15]),
    .local_valid_o         (valid_o[9][15]),
    .local_ready_i         (ready_i[9][15]),
    .credit_upd            (credit_upd)
);

/*Router 9,16*/    
cast_router #(
    .isUBM_list            (isUBM_list_9_16),
    .isFC_list             (isFC_list_9_16),
    .FCdn_list             (FCdn_list_9_16),
    .FCpl_list             (FCpl_list_9_16),
    .rt_file_list          (cast_rt_file_list_9_16)
)router_9_16(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_168_to_169),
    .west_valid_i          (valid_168_to_169),
    .west_ready_o          (ready_169_to_168),
    .west_data_o           (data_169_to_168),
    .west_valid_o          (valid_169_to_168),
    .west_ready_i          (ready_168_to_169),
    .east_data_i           (34'b0),
    .east_valid_i          (1'b0),
    .east_ready_o          (),
    .east_data_o           (),
    .east_valid_o          (),
    .east_ready_i          (1'b0),
    .vert0_data_i          (data_159_to_169_v0),
    .vert0_valid_i         (valid_159_to_169_v0),
    .vert0_ready_o         (ready_169_to_159_v0),
    .vert0_data_o          (data_169_to_179_v0),
    .vert0_valid_o         (valid_169_to_179_v0),
    .vert0_ready_i         (ready_179_to_169_v0),
    .vert1_data_i          (data_159_to_169_v1),
    .vert1_valid_i         (valid_159_to_169_v1),
    .vert1_ready_o         (ready_169_to_159_v1),
    .vert1_data_o          (data_169_to_179_v1),
    .vert1_valid_o         (valid_169_to_179_v1),
    .vert1_ready_i         (ready_179_to_169_v1),
    .local_data_i          (data_i[9][16]),
    .local_valid_i         (valid_i[9][16]),
    .local_ready_o         (ready_o[9][16]),
    .local_data_o          (data_o[9][16]),
    .local_valid_o         (valid_o[9][16]),
    .local_ready_i         (ready_i[9][16]),
    .credit_upd            (credit_upd)
);

/*Router 9,17*/    
cast_router #(
    .isUBM_list            (isUBM_list_9_17),
    .isFC_list             (isFC_list_9_17),
    .FCdn_list             (FCdn_list_9_17),
    .FCpl_list             (FCpl_list_9_17),
    .rt_file_list          (cast_rt_file_list_9_17)
)router_9_17(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_178_to_179),
    .west_valid_i          (valid_178_to_179),
    .west_ready_o          (ready_179_to_178),
    .west_data_o           (data_179_to_178),
    .west_valid_o          (valid_179_to_178),
    .west_ready_i          (ready_178_to_179),
    .east_data_i           (34'b0),
    .east_valid_i          (1'b0),
    .east_ready_o          (),
    .east_data_o           (),
    .east_valid_o          (),
    .east_ready_i          (1'b0),
    .vert0_data_i          (data_169_to_179_v0),
    .vert0_valid_i         (valid_169_to_179_v0),
    .vert0_ready_o         (ready_179_to_169_v0),
    .vert0_data_o          (data_179_to_189_v0),
    .vert0_valid_o         (valid_179_to_189_v0),
    .vert0_ready_i         (ready_189_to_179_v0),
    .vert1_data_i          (data_169_to_179_v1),
    .vert1_valid_i         (valid_169_to_179_v1),
    .vert1_ready_o         (ready_179_to_169_v1),
    .vert1_data_o          (data_179_to_189_v1),
    .vert1_valid_o         (valid_179_to_189_v1),
    .vert1_ready_i         (ready_189_to_179_v1),
    .local_data_i          (data_i[9][17]),
    .local_valid_i         (valid_i[9][17]),
    .local_ready_o         (ready_o[9][17]),
    .local_data_o          (data_o[9][17]),
    .local_valid_o         (valid_o[9][17]),
    .local_ready_i         (ready_i[9][17]),
    .credit_upd            (credit_upd)
);

/*Router 9,18*/    
cast_router #(
    .isUBM_list            (isUBM_list_9_18),
    .isFC_list             (isFC_list_9_18),
    .FCdn_list             (FCdn_list_9_18),
    .FCpl_list             (FCpl_list_9_18),
    .rt_file_list          (cast_rt_file_list_9_18)
)router_9_18(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_188_to_189),
    .west_valid_i          (valid_188_to_189),
    .west_ready_o          (ready_189_to_188),
    .west_data_o           (data_189_to_188),
    .west_valid_o          (valid_189_to_188),
    .west_ready_i          (ready_188_to_189),
    .east_data_i           (34'b0),
    .east_valid_i          (1'b0),
    .east_ready_o          (),
    .east_data_o           (),
    .east_valid_o          (),
    .east_ready_i          (1'b0),
    .vert0_data_i          (data_179_to_189_v0),
    .vert0_valid_i         (valid_179_to_189_v0),
    .vert0_ready_o         (ready_189_to_179_v0),
    .vert0_data_o          (data_189_to_199_v0),
    .vert0_valid_o         (valid_189_to_199_v0),
    .vert0_ready_i         (ready_199_to_189_v0),
    .vert1_data_i          (data_179_to_189_v1),
    .vert1_valid_i         (valid_179_to_189_v1),
    .vert1_ready_o         (ready_189_to_179_v1),
    .vert1_data_o          (data_189_to_199_v1),
    .vert1_valid_o         (valid_189_to_199_v1),
    .vert1_ready_i         (ready_199_to_189_v1),
    .local_data_i          (data_i[9][18]),
    .local_valid_i         (valid_i[9][18]),
    .local_ready_o         (ready_o[9][18]),
    .local_data_o          (data_o[9][18]),
    .local_valid_o         (valid_o[9][18]),
    .local_ready_i         (ready_i[9][18]),
    .credit_upd            (credit_upd)
);

/*Router 9,19*/    
cast_router #(
    .isUBM_list            (isUBM_list_9_19),
    .isFC_list             (isFC_list_9_19),
    .FCdn_list             (FCdn_list_9_19),
    .FCpl_list             (FCpl_list_9_19),
    .rt_file_list          (cast_rt_file_list_9_19)
)router_9_19(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_198_to_199),
    .west_valid_i          (valid_198_to_199),
    .west_ready_o          (ready_199_to_198),
    .west_data_o           (data_199_to_198),
    .west_valid_o          (valid_199_to_198),
    .west_ready_i          (ready_198_to_199),
    .east_data_i           (34'b0),
    .east_valid_i          (1'b0),
    .east_ready_o          (),
    .east_data_o           (),
    .east_valid_o          (),
    .east_ready_i          (1'b0),
    .vert0_data_i          (data_189_to_199_v0),
    .vert0_valid_i         (valid_189_to_199_v0),
    .vert0_ready_o         (ready_199_to_189_v0),
    .vert0_data_o          (data_199_to_209_v0),
    .vert0_valid_o         (valid_199_to_209_v0),
    .vert0_ready_i         (ready_209_to_199_v0),
    .vert1_data_i          (data_189_to_199_v1),
    .vert1_valid_i         (valid_189_to_199_v1),
    .vert1_ready_o         (ready_199_to_189_v1),
    .vert1_data_o          (data_199_to_209_v1),
    .vert1_valid_o         (valid_199_to_209_v1),
    .vert1_ready_i         (ready_209_to_199_v1),
    .local_data_i          (data_i[9][19]),
    .local_valid_i         (valid_i[9][19]),
    .local_ready_o         (ready_o[9][19]),
    .local_data_o          (data_o[9][19]),
    .local_valid_o         (valid_o[9][19]),
    .local_ready_i         (ready_i[9][19]),
    .credit_upd            (credit_upd)
);

/*Router 9,20*/    
cast_router #(
    .isUBM_list            (isUBM_list_9_20),
    .isFC_list             (isFC_list_9_20),
    .FCdn_list             (FCdn_list_9_20),
    .FCpl_list             (FCpl_list_9_20),
    .rt_file_list          (cast_rt_file_list_9_20)
)router_9_20(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_208_to_209),
    .west_valid_i          (valid_208_to_209),
    .west_ready_o          (ready_209_to_208),
    .west_data_o           (data_209_to_208),
    .west_valid_o          (valid_209_to_208),
    .west_ready_i          (ready_208_to_209),
    .east_data_i           (34'b0),
    .east_valid_i          (1'b0),
    .east_ready_o          (),
    .east_data_o           (),
    .east_valid_o          (),
    .east_ready_i          (1'b0),
    .vert0_data_i          (data_199_to_209_v0),
    .vert0_valid_i         (valid_199_to_209_v0),
    .vert0_ready_o         (ready_209_to_199_v0),
    .vert0_data_o          (data_209_to_219_v0),
    .vert0_valid_o         (valid_209_to_219_v0),
    .vert0_ready_i         (ready_219_to_209_v0),
    .vert1_data_i          (data_199_to_209_v1),
    .vert1_valid_i         (valid_199_to_209_v1),
    .vert1_ready_o         (ready_209_to_199_v1),
    .vert1_data_o          (data_209_to_219_v1),
    .vert1_valid_o         (valid_209_to_219_v1),
    .vert1_ready_i         (ready_219_to_209_v1),
    .local_data_i          (data_i[9][20]),
    .local_valid_i         (valid_i[9][20]),
    .local_ready_o         (ready_o[9][20]),
    .local_data_o          (data_o[9][20]),
    .local_valid_o         (valid_o[9][20]),
    .local_ready_i         (ready_i[9][20]),
    .credit_upd            (credit_upd)
);

/*Router 9,21*/    
cast_router #(
    .isUBM_list            (isUBM_list_9_21),
    .isFC_list             (isFC_list_9_21),
    .FCdn_list             (FCdn_list_9_21),
    .FCpl_list             (FCpl_list_9_21),
    .rt_file_list          (cast_rt_file_list_9_21)
)router_9_21(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_218_to_219),
    .west_valid_i          (valid_218_to_219),
    .west_ready_o          (ready_219_to_218),
    .west_data_o           (data_219_to_218),
    .west_valid_o          (valid_219_to_218),
    .west_ready_i          (ready_218_to_219),
    .east_data_i           (34'b0),
    .east_valid_i          (1'b0),
    .east_ready_o          (),
    .east_data_o           (),
    .east_valid_o          (),
    .east_ready_i          (1'b0),
    .vert0_data_i          (data_209_to_219_v0),
    .vert0_valid_i         (valid_209_to_219_v0),
    .vert0_ready_o         (ready_219_to_209_v0),
    .vert0_data_o          (data_219_to_229_v0),
    .vert0_valid_o         (valid_219_to_229_v0),
    .vert0_ready_i         (ready_229_to_219_v0),
    .vert1_data_i          (data_209_to_219_v1),
    .vert1_valid_i         (valid_209_to_219_v1),
    .vert1_ready_o         (ready_219_to_209_v1),
    .vert1_data_o          (data_219_to_229_v1),
    .vert1_valid_o         (valid_219_to_229_v1),
    .vert1_ready_i         (ready_229_to_219_v1),
    .local_data_i          (data_i[9][21]),
    .local_valid_i         (valid_i[9][21]),
    .local_ready_o         (ready_o[9][21]),
    .local_data_o          (data_o[9][21]),
    .local_valid_o         (valid_o[9][21]),
    .local_ready_i         (ready_i[9][21]),
    .credit_upd            (credit_upd)
);

/*Router 9,22*/    
cast_router #(
    .isUBM_list            (isUBM_list_9_22),
    .isFC_list             (isFC_list_9_22),
    .FCdn_list             (FCdn_list_9_22),
    .FCpl_list             (FCpl_list_9_22),
    .rt_file_list          (cast_rt_file_list_9_22)
)router_9_22(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_228_to_229),
    .west_valid_i          (valid_228_to_229),
    .west_ready_o          (ready_229_to_228),
    .west_data_o           (data_o_flee1),
    .west_valid_o          (valid_o_flee1),
    .west_ready_i          (ready_i_flee1),
    .east_data_i           (34'b0),
    .east_valid_i          (1'b0),
    .east_ready_o          (),
    .east_data_o           (),
    .east_valid_o          (),
    .east_ready_i          (1'b0),
    .vert0_data_i          (data_219_to_229_v0),
    .vert0_valid_i         (valid_219_to_229_v0),
    .vert0_ready_o         (ready_229_to_219_v0),
    .vert0_data_o          (data_229_to_239_v0),
    .vert0_valid_o         (valid_229_to_239_v0),
    .vert0_ready_i         (ready_239_to_229_v0),
    .vert1_data_i          (data_219_to_229_v1),
    .vert1_valid_i         (valid_219_to_229_v1),
    .vert1_ready_o         (ready_229_to_219_v1),
    .vert1_data_o          (data_229_to_239_v1),
    .vert1_valid_o         (valid_229_to_239_v1),
    .vert1_ready_i         (ready_239_to_229_v1),
    .local_data_i          (data_i[9][22]),
    .local_valid_i         (valid_i[9][22]),
    .local_ready_o         (ready_o[9][22]),
    .local_data_o          (data_o[9][22]),
    .local_valid_o         (valid_o[9][22]),
    .local_ready_i         (ready_i[9][22]),
    .credit_upd            (credit_upd)
);

/*Router 9,23*/    
cast_router #(
    .isUBM_list            (isUBM_list_9_23),
    .isFC_list             (isFC_list_9_23),
    .FCdn_list             (FCdn_list_9_23),
    .FCpl_list             (FCpl_list_9_23),
    .rt_file_list          (cast_rt_file_list_9_23)
)router_9_23(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_238_to_239),
    .west_valid_i          (valid_238_to_239),
    .west_ready_o          (ready_239_to_238),
    .west_data_o           (data_239_to_238),
    .west_valid_o          (valid_239_to_238),
    .west_ready_i          (ready_238_to_239),
    .east_data_i           (34'b0),
    .east_valid_i          (1'b0),
    .east_ready_o          (),
    .east_data_o           (),
    .east_valid_o          (),
    .east_ready_i          (1'b0),
    .vert0_data_i          (data_229_to_239_v0),
    .vert0_valid_i         (valid_229_to_239_v0),
    .vert0_ready_o         (ready_239_to_229_v0),
    .vert0_data_o          (data_239_to_249_v0),
    .vert0_valid_o         (valid_239_to_249_v0),
    .vert0_ready_i         (ready_249_to_239_v0),
    .vert1_data_i          (data_229_to_239_v1),
    .vert1_valid_i         (valid_229_to_239_v1),
    .vert1_ready_o         (ready_239_to_229_v1),
    .vert1_data_o          (data_239_to_249_v1),
    .vert1_valid_o         (valid_239_to_249_v1),
    .vert1_ready_i         (ready_249_to_239_v1),
    .local_data_i          (data_i[9][23]),
    .local_valid_i         (valid_i[9][23]),
    .local_ready_o         (ready_o[9][23]),
    .local_data_o          (data_o[9][23]),
    .local_valid_o         (valid_o[9][23]),
    .local_ready_i         (ready_i[9][23]),
    .credit_upd            (credit_upd)
);

/*Router 9,24*/    
cast_router #(
    .isUBM_list            (isUBM_list_9_24),
    .isFC_list             (isFC_list_9_24),
    .FCdn_list             (FCdn_list_9_24),
    .FCpl_list             (FCpl_list_9_24),
    .rt_file_list          (cast_rt_file_list_9_24)
)router_9_24(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_248_to_249),
    .west_valid_i          (valid_248_to_249),
    .west_ready_o          (ready_249_to_248),
    .west_data_o           (data_249_to_248),
    .west_valid_o          (valid_249_to_248),
    .west_ready_i          (ready_248_to_249),
    .east_data_i           (34'b0),
    .east_valid_i          (1'b0),
    .east_ready_o          (),
    .east_data_o           (),
    .east_valid_o          (),
    .east_ready_i          (1'b0),
    .vert0_data_i          (data_239_to_249_v0),
    .vert0_valid_i         (valid_239_to_249_v0),
    .vert0_ready_o         (ready_249_to_239_v0),
    .vert0_data_o          (),
    .vert0_valid_o         (),
    .vert0_ready_i         (1'b0),
    .vert1_data_i          (data_239_to_249_v1),
    .vert1_valid_i         (valid_239_to_249_v1),
    .vert1_ready_o         (ready_249_to_239_v1),
    .vert1_data_o          (),
    .vert1_valid_o         (),
    .vert1_ready_i         (1'b0),
    .local_data_i          (data_i[9][24]),
    .local_valid_i         (valid_i[9][24]),
    .local_ready_o         (ready_o[9][24]),
    .local_data_o          (data_o[9][24]),
    .local_valid_o         (valid_o[9][24]),
    .local_ready_i         (ready_i[9][24]),
    .credit_upd            (credit_upd)
);

endmodule
