`include "params.svh"
`include "network_config.svh"

module system (
    input       wire                            clk,
    input       wire                            rstn,

    input       wire        [`DW-1:0]           data_i_stab,
    input       wire                            valid_i_stab,
    output      wire                            ready_o_stab,

    output      wire        [`DW-1:0]           data_o_flee0,
    output      wire                            valid_o_flee0,
    input       wire                            ready_i_flee0,
    output      wire        [`DW-1:0]           data_o_flee1,
    output      wire                            valid_o_flee1,
    input       wire                            ready_i_flee1,
    output      wire        [`DW-1:0]           data_o_flee2,
    output      wire                            valid_o_flee2,
    input       wire                            ready_i_flee2,
    output      wire        [`DW-1:0]           data_o_flee3,
    output      wire                            valid_o_flee3,
    input       wire                            ready_i_flee3,
    output      wire        [`DW-1:0]           data_o_flee4,
    output      wire                            valid_o_flee4,
    input       wire                            ready_i_flee4,
    output      wire        [`DW-1:0]           data_o_flee5,
    output      wire                            valid_o_flee5,
    input       wire                            ready_i_flee5,
    output      wire        [`DW-1:0]           data_o_flee6,
    output      wire                            valid_o_flee6,
    input       wire                            ready_i_flee6,
    output      wire        [`DW-1:0]           data_o_flee7,
    output      wire                            valid_o_flee7,
    input       wire                            ready_i_flee7
);

wire [`DW-1:0] cast_data_pe_2_nw[`NOC_WIDTH][`NOC_HEIGHT], merge_data_pe_2_nw[`NOC_WIDTH][`NOC_HEIGHT], gather_data_pe_2_nw[`NOC_WIDTH][`NOC_HEIGHT], cast_data_nw_2_pe[`NOC_WIDTH][`NOC_HEIGHT], merge_data_nw_2_pe[`NOC_WIDTH][`NOC_HEIGHT], gather_data_nw_2_pe[`NOC_WIDTH][`NOC_HEIGHT];
wire  cast_valid_pe_2_nw[`NOC_WIDTH][`NOC_HEIGHT], merge_valid_pe_2_nw[`NOC_WIDTH][`NOC_HEIGHT], gather_valid_pe_2_nw[`NOC_WIDTH][`NOC_HEIGHT], cast_valid_nw_2_pe[`NOC_WIDTH][`NOC_HEIGHT], merge_valid_nw_2_pe[`NOC_WIDTH][`NOC_HEIGHT], gather_valid_nw_2_pe[`NOC_WIDTH][`NOC_HEIGHT];
wire  cast_ready_pe_2_nw[`NOC_WIDTH][`NOC_HEIGHT], merge_ready_pe_2_nw[`NOC_WIDTH][`NOC_HEIGHT], gather_ready_pe_2_nw[`NOC_WIDTH][`NOC_HEIGHT], cast_ready_nw_2_pe[`NOC_WIDTH][`NOC_HEIGHT], merge_ready_nw_2_pe[`NOC_WIDTH][`NOC_HEIGHT], gather_ready_nw_2_pe[`NOC_WIDTH][`NOC_HEIGHT];

network nw(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .data_i_stab                                       (data_i_stab),
    .valid_i_stab                                      (valid_i_stab),
    .ready_o_stab                                      (ready_o_stab),
    .data_o_flee0                                      (data_o_flee0),
    .valid_o_flee0                                     (valid_o_flee0),
    .ready_i_flee0                                     (ready_i_flee0),
    .data_o_flee1                                      (data_o_flee1),
    .valid_o_flee1                                     (valid_o_flee1),
    .ready_i_flee1                                     (ready_i_flee1),
    .data_o_flee2                                      (data_o_flee2),
    .valid_o_flee2                                     (valid_o_flee2),
    .ready_i_flee2                                     (ready_i_flee2),
    .data_o_flee3                                      (data_o_flee3),
    .valid_o_flee3                                     (valid_o_flee3),
    .ready_i_flee3                                     (ready_i_flee3),
    .data_o_flee4                                      (data_o_flee4),
    .valid_o_flee4                                     (valid_o_flee4),
    .ready_i_flee4                                     (ready_i_flee4),
    .data_o_flee5                                      (data_o_flee5),
    .valid_o_flee5                                     (valid_o_flee5),
    .ready_i_flee5                                     (ready_i_flee5),
    .data_o_flee6                                      (data_o_flee6),
    .valid_o_flee6                                     (valid_o_flee6),
    .ready_i_flee6                                     (ready_i_flee6),
    .data_o_flee7                                      (data_o_flee7),
    .valid_o_flee7                                     (valid_o_flee7),
    .ready_i_flee7                                     (ready_i_flee7),
    .cast_data_i_0_0                               (cast_data_pe_2_nw[0][0]),
    .cast_valid_i_0_0                              (cast_valid_pe_2_nw[0][0]),
    .cast_ready_o_0_0                              (cast_ready_nw_2_pe[0][0]),
    .merge_data_i_0_0                              (merge_data_pe_2_nw[0][0]),
    .merge_valid_i_0_0                             (merge_valid_pe_2_nw[0][0]),
    .merge_ready_o_0_0                             (merge_ready_nw_2_pe[0][0]),
    .gather_data_i_0_0                             (gather_data_pe_2_nw[0][0]),
    .gather_valid_i_0_0                            (gather_valid_pe_2_nw[0][0]),
    .gather_ready_o_0_0                            (gather_ready_nw_2_pe[0][0]),

    .cast_data_o_0_0                               (cast_data_nw_2_pe[0][0]),
    .cast_valid_o_0_0                              (cast_valid_nw_2_pe[0][0]),
    .cast_ready_i_0_0                              (cast_ready_pe_2_nw[0][0]),
    .merge_data_o_0_0                              (merge_data_nw_2_pe[0][0]),
    .merge_valid_o_0_0                             (merge_valid_nw_2_pe[0][0]),
    .merge_ready_i_0_0                             (merge_ready_pe_2_nw[0][0]),
    .gather_data_o_0_0                             (gather_data_nw_2_pe[0][0]),
    .gather_valid_o_0_0                            (gather_valid_nw_2_pe[0][0]),
    .gather_ready_i_0_0                            (gather_ready_pe_2_nw[0][0]),
    .cast_data_i_0_1                               (cast_data_pe_2_nw[0][1]),
    .cast_valid_i_0_1                              (cast_valid_pe_2_nw[0][1]),
    .cast_ready_o_0_1                              (cast_ready_nw_2_pe[0][1]),
    .merge_data_i_0_1                              (merge_data_pe_2_nw[0][1]),
    .merge_valid_i_0_1                             (merge_valid_pe_2_nw[0][1]),
    .merge_ready_o_0_1                             (merge_ready_nw_2_pe[0][1]),
    .gather_data_i_0_1                             (gather_data_pe_2_nw[0][1]),
    .gather_valid_i_0_1                            (gather_valid_pe_2_nw[0][1]),
    .gather_ready_o_0_1                            (gather_ready_nw_2_pe[0][1]),

    .cast_data_o_0_1                               (cast_data_nw_2_pe[0][1]),
    .cast_valid_o_0_1                              (cast_valid_nw_2_pe[0][1]),
    .cast_ready_i_0_1                              (cast_ready_pe_2_nw[0][1]),
    .merge_data_o_0_1                              (merge_data_nw_2_pe[0][1]),
    .merge_valid_o_0_1                             (merge_valid_nw_2_pe[0][1]),
    .merge_ready_i_0_1                             (merge_ready_pe_2_nw[0][1]),
    .gather_data_o_0_1                             (gather_data_nw_2_pe[0][1]),
    .gather_valid_o_0_1                            (gather_valid_nw_2_pe[0][1]),
    .gather_ready_i_0_1                            (gather_ready_pe_2_nw[0][1]),
    .cast_data_i_0_2                               (cast_data_pe_2_nw[0][2]),
    .cast_valid_i_0_2                              (cast_valid_pe_2_nw[0][2]),
    .cast_ready_o_0_2                              (cast_ready_nw_2_pe[0][2]),
    .merge_data_i_0_2                              (merge_data_pe_2_nw[0][2]),
    .merge_valid_i_0_2                             (merge_valid_pe_2_nw[0][2]),
    .merge_ready_o_0_2                             (merge_ready_nw_2_pe[0][2]),
    .gather_data_i_0_2                             (gather_data_pe_2_nw[0][2]),
    .gather_valid_i_0_2                            (gather_valid_pe_2_nw[0][2]),
    .gather_ready_o_0_2                            (gather_ready_nw_2_pe[0][2]),

    .cast_data_o_0_2                               (cast_data_nw_2_pe[0][2]),
    .cast_valid_o_0_2                              (cast_valid_nw_2_pe[0][2]),
    .cast_ready_i_0_2                              (cast_ready_pe_2_nw[0][2]),
    .merge_data_o_0_2                              (merge_data_nw_2_pe[0][2]),
    .merge_valid_o_0_2                             (merge_valid_nw_2_pe[0][2]),
    .merge_ready_i_0_2                             (merge_ready_pe_2_nw[0][2]),
    .gather_data_o_0_2                             (gather_data_nw_2_pe[0][2]),
    .gather_valid_o_0_2                            (gather_valid_nw_2_pe[0][2]),
    .gather_ready_i_0_2                            (gather_ready_pe_2_nw[0][2]),
    .cast_data_i_0_3                               (cast_data_pe_2_nw[0][3]),
    .cast_valid_i_0_3                              (cast_valid_pe_2_nw[0][3]),
    .cast_ready_o_0_3                              (cast_ready_nw_2_pe[0][3]),
    .merge_data_i_0_3                              (merge_data_pe_2_nw[0][3]),
    .merge_valid_i_0_3                             (merge_valid_pe_2_nw[0][3]),
    .merge_ready_o_0_3                             (merge_ready_nw_2_pe[0][3]),
    .gather_data_i_0_3                             (gather_data_pe_2_nw[0][3]),
    .gather_valid_i_0_3                            (gather_valid_pe_2_nw[0][3]),
    .gather_ready_o_0_3                            (gather_ready_nw_2_pe[0][3]),

    .cast_data_o_0_3                               (cast_data_nw_2_pe[0][3]),
    .cast_valid_o_0_3                              (cast_valid_nw_2_pe[0][3]),
    .cast_ready_i_0_3                              (cast_ready_pe_2_nw[0][3]),
    .merge_data_o_0_3                              (merge_data_nw_2_pe[0][3]),
    .merge_valid_o_0_3                             (merge_valid_nw_2_pe[0][3]),
    .merge_ready_i_0_3                             (merge_ready_pe_2_nw[0][3]),
    .gather_data_o_0_3                             (gather_data_nw_2_pe[0][3]),
    .gather_valid_o_0_3                            (gather_valid_nw_2_pe[0][3]),
    .gather_ready_i_0_3                            (gather_ready_pe_2_nw[0][3]),
    .cast_data_i_0_4                               (cast_data_pe_2_nw[0][4]),
    .cast_valid_i_0_4                              (cast_valid_pe_2_nw[0][4]),
    .cast_ready_o_0_4                              (cast_ready_nw_2_pe[0][4]),
    .merge_data_i_0_4                              (merge_data_pe_2_nw[0][4]),
    .merge_valid_i_0_4                             (merge_valid_pe_2_nw[0][4]),
    .merge_ready_o_0_4                             (merge_ready_nw_2_pe[0][4]),
    .gather_data_i_0_4                             (gather_data_pe_2_nw[0][4]),
    .gather_valid_i_0_4                            (gather_valid_pe_2_nw[0][4]),
    .gather_ready_o_0_4                            (gather_ready_nw_2_pe[0][4]),

    .cast_data_o_0_4                               (cast_data_nw_2_pe[0][4]),
    .cast_valid_o_0_4                              (cast_valid_nw_2_pe[0][4]),
    .cast_ready_i_0_4                              (cast_ready_pe_2_nw[0][4]),
    .merge_data_o_0_4                              (merge_data_nw_2_pe[0][4]),
    .merge_valid_o_0_4                             (merge_valid_nw_2_pe[0][4]),
    .merge_ready_i_0_4                             (merge_ready_pe_2_nw[0][4]),
    .gather_data_o_0_4                             (gather_data_nw_2_pe[0][4]),
    .gather_valid_o_0_4                            (gather_valid_nw_2_pe[0][4]),
    .gather_ready_i_0_4                            (gather_ready_pe_2_nw[0][4]),
    .cast_data_i_0_5                               (cast_data_pe_2_nw[0][5]),
    .cast_valid_i_0_5                              (cast_valid_pe_2_nw[0][5]),
    .cast_ready_o_0_5                              (cast_ready_nw_2_pe[0][5]),
    .merge_data_i_0_5                              (merge_data_pe_2_nw[0][5]),
    .merge_valid_i_0_5                             (merge_valid_pe_2_nw[0][5]),
    .merge_ready_o_0_5                             (merge_ready_nw_2_pe[0][5]),
    .gather_data_i_0_5                             (gather_data_pe_2_nw[0][5]),
    .gather_valid_i_0_5                            (gather_valid_pe_2_nw[0][5]),
    .gather_ready_o_0_5                            (gather_ready_nw_2_pe[0][5]),

    .cast_data_o_0_5                               (cast_data_nw_2_pe[0][5]),
    .cast_valid_o_0_5                              (cast_valid_nw_2_pe[0][5]),
    .cast_ready_i_0_5                              (cast_ready_pe_2_nw[0][5]),
    .merge_data_o_0_5                              (merge_data_nw_2_pe[0][5]),
    .merge_valid_o_0_5                             (merge_valid_nw_2_pe[0][5]),
    .merge_ready_i_0_5                             (merge_ready_pe_2_nw[0][5]),
    .gather_data_o_0_5                             (gather_data_nw_2_pe[0][5]),
    .gather_valid_o_0_5                            (gather_valid_nw_2_pe[0][5]),
    .gather_ready_i_0_5                            (gather_ready_pe_2_nw[0][5]),
    .cast_data_i_0_6                               (cast_data_pe_2_nw[0][6]),
    .cast_valid_i_0_6                              (cast_valid_pe_2_nw[0][6]),
    .cast_ready_o_0_6                              (cast_ready_nw_2_pe[0][6]),
    .merge_data_i_0_6                              (merge_data_pe_2_nw[0][6]),
    .merge_valid_i_0_6                             (merge_valid_pe_2_nw[0][6]),
    .merge_ready_o_0_6                             (merge_ready_nw_2_pe[0][6]),
    .gather_data_i_0_6                             (gather_data_pe_2_nw[0][6]),
    .gather_valid_i_0_6                            (gather_valid_pe_2_nw[0][6]),
    .gather_ready_o_0_6                            (gather_ready_nw_2_pe[0][6]),

    .cast_data_o_0_6                               (cast_data_nw_2_pe[0][6]),
    .cast_valid_o_0_6                              (cast_valid_nw_2_pe[0][6]),
    .cast_ready_i_0_6                              (cast_ready_pe_2_nw[0][6]),
    .merge_data_o_0_6                              (merge_data_nw_2_pe[0][6]),
    .merge_valid_o_0_6                             (merge_valid_nw_2_pe[0][6]),
    .merge_ready_i_0_6                             (merge_ready_pe_2_nw[0][6]),
    .gather_data_o_0_6                             (gather_data_nw_2_pe[0][6]),
    .gather_valid_o_0_6                            (gather_valid_nw_2_pe[0][6]),
    .gather_ready_i_0_6                            (gather_ready_pe_2_nw[0][6]),
    .cast_data_i_0_7                               (cast_data_pe_2_nw[0][7]),
    .cast_valid_i_0_7                              (cast_valid_pe_2_nw[0][7]),
    .cast_ready_o_0_7                              (cast_ready_nw_2_pe[0][7]),
    .merge_data_i_0_7                              (merge_data_pe_2_nw[0][7]),
    .merge_valid_i_0_7                             (merge_valid_pe_2_nw[0][7]),
    .merge_ready_o_0_7                             (merge_ready_nw_2_pe[0][7]),
    .gather_data_i_0_7                             (gather_data_pe_2_nw[0][7]),
    .gather_valid_i_0_7                            (gather_valid_pe_2_nw[0][7]),
    .gather_ready_o_0_7                            (gather_ready_nw_2_pe[0][7]),

    .cast_data_o_0_7                               (cast_data_nw_2_pe[0][7]),
    .cast_valid_o_0_7                              (cast_valid_nw_2_pe[0][7]),
    .cast_ready_i_0_7                              (cast_ready_pe_2_nw[0][7]),
    .merge_data_o_0_7                              (merge_data_nw_2_pe[0][7]),
    .merge_valid_o_0_7                             (merge_valid_nw_2_pe[0][7]),
    .merge_ready_i_0_7                             (merge_ready_pe_2_nw[0][7]),
    .gather_data_o_0_7                             (gather_data_nw_2_pe[0][7]),
    .gather_valid_o_0_7                            (gather_valid_nw_2_pe[0][7]),
    .gather_ready_i_0_7                            (gather_ready_pe_2_nw[0][7]),
    .cast_data_i_0_8                               (cast_data_pe_2_nw[0][8]),
    .cast_valid_i_0_8                              (cast_valid_pe_2_nw[0][8]),
    .cast_ready_o_0_8                              (cast_ready_nw_2_pe[0][8]),
    .merge_data_i_0_8                              (merge_data_pe_2_nw[0][8]),
    .merge_valid_i_0_8                             (merge_valid_pe_2_nw[0][8]),
    .merge_ready_o_0_8                             (merge_ready_nw_2_pe[0][8]),
    .gather_data_i_0_8                             (gather_data_pe_2_nw[0][8]),
    .gather_valid_i_0_8                            (gather_valid_pe_2_nw[0][8]),
    .gather_ready_o_0_8                            (gather_ready_nw_2_pe[0][8]),

    .cast_data_o_0_8                               (cast_data_nw_2_pe[0][8]),
    .cast_valid_o_0_8                              (cast_valid_nw_2_pe[0][8]),
    .cast_ready_i_0_8                              (cast_ready_pe_2_nw[0][8]),
    .merge_data_o_0_8                              (merge_data_nw_2_pe[0][8]),
    .merge_valid_o_0_8                             (merge_valid_nw_2_pe[0][8]),
    .merge_ready_i_0_8                             (merge_ready_pe_2_nw[0][8]),
    .gather_data_o_0_8                             (gather_data_nw_2_pe[0][8]),
    .gather_valid_o_0_8                            (gather_valid_nw_2_pe[0][8]),
    .gather_ready_i_0_8                            (gather_ready_pe_2_nw[0][8]),
    .cast_data_i_0_9                               (cast_data_pe_2_nw[0][9]),
    .cast_valid_i_0_9                              (cast_valid_pe_2_nw[0][9]),
    .cast_ready_o_0_9                              (cast_ready_nw_2_pe[0][9]),
    .merge_data_i_0_9                              (merge_data_pe_2_nw[0][9]),
    .merge_valid_i_0_9                             (merge_valid_pe_2_nw[0][9]),
    .merge_ready_o_0_9                             (merge_ready_nw_2_pe[0][9]),
    .gather_data_i_0_9                             (gather_data_pe_2_nw[0][9]),
    .gather_valid_i_0_9                            (gather_valid_pe_2_nw[0][9]),
    .gather_ready_o_0_9                            (gather_ready_nw_2_pe[0][9]),

    .cast_data_o_0_9                               (cast_data_nw_2_pe[0][9]),
    .cast_valid_o_0_9                              (cast_valid_nw_2_pe[0][9]),
    .cast_ready_i_0_9                              (cast_ready_pe_2_nw[0][9]),
    .merge_data_o_0_9                              (merge_data_nw_2_pe[0][9]),
    .merge_valid_o_0_9                             (merge_valid_nw_2_pe[0][9]),
    .merge_ready_i_0_9                             (merge_ready_pe_2_nw[0][9]),
    .gather_data_o_0_9                             (gather_data_nw_2_pe[0][9]),
    .gather_valid_o_0_9                            (gather_valid_nw_2_pe[0][9]),
    .gather_ready_i_0_9                            (gather_ready_pe_2_nw[0][9]),
    .cast_data_i_0_10                               (cast_data_pe_2_nw[0][10]),
    .cast_valid_i_0_10                              (cast_valid_pe_2_nw[0][10]),
    .cast_ready_o_0_10                              (cast_ready_nw_2_pe[0][10]),
    .merge_data_i_0_10                              (merge_data_pe_2_nw[0][10]),
    .merge_valid_i_0_10                             (merge_valid_pe_2_nw[0][10]),
    .merge_ready_o_0_10                             (merge_ready_nw_2_pe[0][10]),
    .gather_data_i_0_10                             (gather_data_pe_2_nw[0][10]),
    .gather_valid_i_0_10                            (gather_valid_pe_2_nw[0][10]),
    .gather_ready_o_0_10                            (gather_ready_nw_2_pe[0][10]),

    .cast_data_o_0_10                               (cast_data_nw_2_pe[0][10]),
    .cast_valid_o_0_10                              (cast_valid_nw_2_pe[0][10]),
    .cast_ready_i_0_10                              (cast_ready_pe_2_nw[0][10]),
    .merge_data_o_0_10                              (merge_data_nw_2_pe[0][10]),
    .merge_valid_o_0_10                             (merge_valid_nw_2_pe[0][10]),
    .merge_ready_i_0_10                             (merge_ready_pe_2_nw[0][10]),
    .gather_data_o_0_10                             (gather_data_nw_2_pe[0][10]),
    .gather_valid_o_0_10                            (gather_valid_nw_2_pe[0][10]),
    .gather_ready_i_0_10                            (gather_ready_pe_2_nw[0][10]),
    .cast_data_i_0_11                               (cast_data_pe_2_nw[0][11]),
    .cast_valid_i_0_11                              (cast_valid_pe_2_nw[0][11]),
    .cast_ready_o_0_11                              (cast_ready_nw_2_pe[0][11]),
    .merge_data_i_0_11                              (merge_data_pe_2_nw[0][11]),
    .merge_valid_i_0_11                             (merge_valid_pe_2_nw[0][11]),
    .merge_ready_o_0_11                             (merge_ready_nw_2_pe[0][11]),
    .gather_data_i_0_11                             (gather_data_pe_2_nw[0][11]),
    .gather_valid_i_0_11                            (gather_valid_pe_2_nw[0][11]),
    .gather_ready_o_0_11                            (gather_ready_nw_2_pe[0][11]),

    .cast_data_o_0_11                               (cast_data_nw_2_pe[0][11]),
    .cast_valid_o_0_11                              (cast_valid_nw_2_pe[0][11]),
    .cast_ready_i_0_11                              (cast_ready_pe_2_nw[0][11]),
    .merge_data_o_0_11                              (merge_data_nw_2_pe[0][11]),
    .merge_valid_o_0_11                             (merge_valid_nw_2_pe[0][11]),
    .merge_ready_i_0_11                             (merge_ready_pe_2_nw[0][11]),
    .gather_data_o_0_11                             (gather_data_nw_2_pe[0][11]),
    .gather_valid_o_0_11                            (gather_valid_nw_2_pe[0][11]),
    .gather_ready_i_0_11                            (gather_ready_pe_2_nw[0][11]),
    .cast_data_i_0_12                               (cast_data_pe_2_nw[0][12]),
    .cast_valid_i_0_12                              (cast_valid_pe_2_nw[0][12]),
    .cast_ready_o_0_12                              (cast_ready_nw_2_pe[0][12]),
    .merge_data_i_0_12                              (merge_data_pe_2_nw[0][12]),
    .merge_valid_i_0_12                             (merge_valid_pe_2_nw[0][12]),
    .merge_ready_o_0_12                             (merge_ready_nw_2_pe[0][12]),
    .gather_data_i_0_12                             (gather_data_pe_2_nw[0][12]),
    .gather_valid_i_0_12                            (gather_valid_pe_2_nw[0][12]),
    .gather_ready_o_0_12                            (gather_ready_nw_2_pe[0][12]),

    .cast_data_o_0_12                               (cast_data_nw_2_pe[0][12]),
    .cast_valid_o_0_12                              (cast_valid_nw_2_pe[0][12]),
    .cast_ready_i_0_12                              (cast_ready_pe_2_nw[0][12]),
    .merge_data_o_0_12                              (merge_data_nw_2_pe[0][12]),
    .merge_valid_o_0_12                             (merge_valid_nw_2_pe[0][12]),
    .merge_ready_i_0_12                             (merge_ready_pe_2_nw[0][12]),
    .gather_data_o_0_12                             (gather_data_nw_2_pe[0][12]),
    .gather_valid_o_0_12                            (gather_valid_nw_2_pe[0][12]),
    .gather_ready_i_0_12                            (gather_ready_pe_2_nw[0][12]),
    .cast_data_i_0_13                               (cast_data_pe_2_nw[0][13]),
    .cast_valid_i_0_13                              (cast_valid_pe_2_nw[0][13]),
    .cast_ready_o_0_13                              (cast_ready_nw_2_pe[0][13]),
    .merge_data_i_0_13                              (merge_data_pe_2_nw[0][13]),
    .merge_valid_i_0_13                             (merge_valid_pe_2_nw[0][13]),
    .merge_ready_o_0_13                             (merge_ready_nw_2_pe[0][13]),
    .gather_data_i_0_13                             (gather_data_pe_2_nw[0][13]),
    .gather_valid_i_0_13                            (gather_valid_pe_2_nw[0][13]),
    .gather_ready_o_0_13                            (gather_ready_nw_2_pe[0][13]),

    .cast_data_o_0_13                               (cast_data_nw_2_pe[0][13]),
    .cast_valid_o_0_13                              (cast_valid_nw_2_pe[0][13]),
    .cast_ready_i_0_13                              (cast_ready_pe_2_nw[0][13]),
    .merge_data_o_0_13                              (merge_data_nw_2_pe[0][13]),
    .merge_valid_o_0_13                             (merge_valid_nw_2_pe[0][13]),
    .merge_ready_i_0_13                             (merge_ready_pe_2_nw[0][13]),
    .gather_data_o_0_13                             (gather_data_nw_2_pe[0][13]),
    .gather_valid_o_0_13                            (gather_valid_nw_2_pe[0][13]),
    .gather_ready_i_0_13                            (gather_ready_pe_2_nw[0][13]),
    .cast_data_i_0_14                               (cast_data_pe_2_nw[0][14]),
    .cast_valid_i_0_14                              (cast_valid_pe_2_nw[0][14]),
    .cast_ready_o_0_14                              (cast_ready_nw_2_pe[0][14]),
    .merge_data_i_0_14                              (merge_data_pe_2_nw[0][14]),
    .merge_valid_i_0_14                             (merge_valid_pe_2_nw[0][14]),
    .merge_ready_o_0_14                             (merge_ready_nw_2_pe[0][14]),
    .gather_data_i_0_14                             (gather_data_pe_2_nw[0][14]),
    .gather_valid_i_0_14                            (gather_valid_pe_2_nw[0][14]),
    .gather_ready_o_0_14                            (gather_ready_nw_2_pe[0][14]),

    .cast_data_o_0_14                               (cast_data_nw_2_pe[0][14]),
    .cast_valid_o_0_14                              (cast_valid_nw_2_pe[0][14]),
    .cast_ready_i_0_14                              (cast_ready_pe_2_nw[0][14]),
    .merge_data_o_0_14                              (merge_data_nw_2_pe[0][14]),
    .merge_valid_o_0_14                             (merge_valid_nw_2_pe[0][14]),
    .merge_ready_i_0_14                             (merge_ready_pe_2_nw[0][14]),
    .gather_data_o_0_14                             (gather_data_nw_2_pe[0][14]),
    .gather_valid_o_0_14                            (gather_valid_nw_2_pe[0][14]),
    .gather_ready_i_0_14                            (gather_ready_pe_2_nw[0][14]),
    .cast_data_i_0_15                               (cast_data_pe_2_nw[0][15]),
    .cast_valid_i_0_15                              (cast_valid_pe_2_nw[0][15]),
    .cast_ready_o_0_15                              (cast_ready_nw_2_pe[0][15]),
    .merge_data_i_0_15                              (merge_data_pe_2_nw[0][15]),
    .merge_valid_i_0_15                             (merge_valid_pe_2_nw[0][15]),
    .merge_ready_o_0_15                             (merge_ready_nw_2_pe[0][15]),
    .gather_data_i_0_15                             (gather_data_pe_2_nw[0][15]),
    .gather_valid_i_0_15                            (gather_valid_pe_2_nw[0][15]),
    .gather_ready_o_0_15                            (gather_ready_nw_2_pe[0][15]),

    .cast_data_o_0_15                               (cast_data_nw_2_pe[0][15]),
    .cast_valid_o_0_15                              (cast_valid_nw_2_pe[0][15]),
    .cast_ready_i_0_15                              (cast_ready_pe_2_nw[0][15]),
    .merge_data_o_0_15                              (merge_data_nw_2_pe[0][15]),
    .merge_valid_o_0_15                             (merge_valid_nw_2_pe[0][15]),
    .merge_ready_i_0_15                             (merge_ready_pe_2_nw[0][15]),
    .gather_data_o_0_15                             (gather_data_nw_2_pe[0][15]),
    .gather_valid_o_0_15                            (gather_valid_nw_2_pe[0][15]),
    .gather_ready_i_0_15                            (gather_ready_pe_2_nw[0][15]),
    .cast_data_i_0_16                               (cast_data_pe_2_nw[0][16]),
    .cast_valid_i_0_16                              (cast_valid_pe_2_nw[0][16]),
    .cast_ready_o_0_16                              (cast_ready_nw_2_pe[0][16]),
    .merge_data_i_0_16                              (merge_data_pe_2_nw[0][16]),
    .merge_valid_i_0_16                             (merge_valid_pe_2_nw[0][16]),
    .merge_ready_o_0_16                             (merge_ready_nw_2_pe[0][16]),
    .gather_data_i_0_16                             (gather_data_pe_2_nw[0][16]),
    .gather_valid_i_0_16                            (gather_valid_pe_2_nw[0][16]),
    .gather_ready_o_0_16                            (gather_ready_nw_2_pe[0][16]),

    .cast_data_o_0_16                               (cast_data_nw_2_pe[0][16]),
    .cast_valid_o_0_16                              (cast_valid_nw_2_pe[0][16]),
    .cast_ready_i_0_16                              (cast_ready_pe_2_nw[0][16]),
    .merge_data_o_0_16                              (merge_data_nw_2_pe[0][16]),
    .merge_valid_o_0_16                             (merge_valid_nw_2_pe[0][16]),
    .merge_ready_i_0_16                             (merge_ready_pe_2_nw[0][16]),
    .gather_data_o_0_16                             (gather_data_nw_2_pe[0][16]),
    .gather_valid_o_0_16                            (gather_valid_nw_2_pe[0][16]),
    .gather_ready_i_0_16                            (gather_ready_pe_2_nw[0][16]),
    .cast_data_i_0_17                               (cast_data_pe_2_nw[0][17]),
    .cast_valid_i_0_17                              (cast_valid_pe_2_nw[0][17]),
    .cast_ready_o_0_17                              (cast_ready_nw_2_pe[0][17]),
    .merge_data_i_0_17                              (merge_data_pe_2_nw[0][17]),
    .merge_valid_i_0_17                             (merge_valid_pe_2_nw[0][17]),
    .merge_ready_o_0_17                             (merge_ready_nw_2_pe[0][17]),
    .gather_data_i_0_17                             (gather_data_pe_2_nw[0][17]),
    .gather_valid_i_0_17                            (gather_valid_pe_2_nw[0][17]),
    .gather_ready_o_0_17                            (gather_ready_nw_2_pe[0][17]),

    .cast_data_o_0_17                               (cast_data_nw_2_pe[0][17]),
    .cast_valid_o_0_17                              (cast_valid_nw_2_pe[0][17]),
    .cast_ready_i_0_17                              (cast_ready_pe_2_nw[0][17]),
    .merge_data_o_0_17                              (merge_data_nw_2_pe[0][17]),
    .merge_valid_o_0_17                             (merge_valid_nw_2_pe[0][17]),
    .merge_ready_i_0_17                             (merge_ready_pe_2_nw[0][17]),
    .gather_data_o_0_17                             (gather_data_nw_2_pe[0][17]),
    .gather_valid_o_0_17                            (gather_valid_nw_2_pe[0][17]),
    .gather_ready_i_0_17                            (gather_ready_pe_2_nw[0][17]),
    .cast_data_i_0_18                               (cast_data_pe_2_nw[0][18]),
    .cast_valid_i_0_18                              (cast_valid_pe_2_nw[0][18]),
    .cast_ready_o_0_18                              (cast_ready_nw_2_pe[0][18]),
    .merge_data_i_0_18                              (merge_data_pe_2_nw[0][18]),
    .merge_valid_i_0_18                             (merge_valid_pe_2_nw[0][18]),
    .merge_ready_o_0_18                             (merge_ready_nw_2_pe[0][18]),
    .gather_data_i_0_18                             (gather_data_pe_2_nw[0][18]),
    .gather_valid_i_0_18                            (gather_valid_pe_2_nw[0][18]),
    .gather_ready_o_0_18                            (gather_ready_nw_2_pe[0][18]),

    .cast_data_o_0_18                               (cast_data_nw_2_pe[0][18]),
    .cast_valid_o_0_18                              (cast_valid_nw_2_pe[0][18]),
    .cast_ready_i_0_18                              (cast_ready_pe_2_nw[0][18]),
    .merge_data_o_0_18                              (merge_data_nw_2_pe[0][18]),
    .merge_valid_o_0_18                             (merge_valid_nw_2_pe[0][18]),
    .merge_ready_i_0_18                             (merge_ready_pe_2_nw[0][18]),
    .gather_data_o_0_18                             (gather_data_nw_2_pe[0][18]),
    .gather_valid_o_0_18                            (gather_valid_nw_2_pe[0][18]),
    .gather_ready_i_0_18                            (gather_ready_pe_2_nw[0][18]),
    .cast_data_i_0_19                               (cast_data_pe_2_nw[0][19]),
    .cast_valid_i_0_19                              (cast_valid_pe_2_nw[0][19]),
    .cast_ready_o_0_19                              (cast_ready_nw_2_pe[0][19]),
    .merge_data_i_0_19                              (merge_data_pe_2_nw[0][19]),
    .merge_valid_i_0_19                             (merge_valid_pe_2_nw[0][19]),
    .merge_ready_o_0_19                             (merge_ready_nw_2_pe[0][19]),
    .gather_data_i_0_19                             (gather_data_pe_2_nw[0][19]),
    .gather_valid_i_0_19                            (gather_valid_pe_2_nw[0][19]),
    .gather_ready_o_0_19                            (gather_ready_nw_2_pe[0][19]),

    .cast_data_o_0_19                               (cast_data_nw_2_pe[0][19]),
    .cast_valid_o_0_19                              (cast_valid_nw_2_pe[0][19]),
    .cast_ready_i_0_19                              (cast_ready_pe_2_nw[0][19]),
    .merge_data_o_0_19                              (merge_data_nw_2_pe[0][19]),
    .merge_valid_o_0_19                             (merge_valid_nw_2_pe[0][19]),
    .merge_ready_i_0_19                             (merge_ready_pe_2_nw[0][19]),
    .gather_data_o_0_19                             (gather_data_nw_2_pe[0][19]),
    .gather_valid_o_0_19                            (gather_valid_nw_2_pe[0][19]),
    .gather_ready_i_0_19                            (gather_ready_pe_2_nw[0][19]),
    .cast_data_i_0_20                               (cast_data_pe_2_nw[0][20]),
    .cast_valid_i_0_20                              (cast_valid_pe_2_nw[0][20]),
    .cast_ready_o_0_20                              (cast_ready_nw_2_pe[0][20]),
    .merge_data_i_0_20                              (merge_data_pe_2_nw[0][20]),
    .merge_valid_i_0_20                             (merge_valid_pe_2_nw[0][20]),
    .merge_ready_o_0_20                             (merge_ready_nw_2_pe[0][20]),
    .gather_data_i_0_20                             (gather_data_pe_2_nw[0][20]),
    .gather_valid_i_0_20                            (gather_valid_pe_2_nw[0][20]),
    .gather_ready_o_0_20                            (gather_ready_nw_2_pe[0][20]),

    .cast_data_o_0_20                               (cast_data_nw_2_pe[0][20]),
    .cast_valid_o_0_20                              (cast_valid_nw_2_pe[0][20]),
    .cast_ready_i_0_20                              (cast_ready_pe_2_nw[0][20]),
    .merge_data_o_0_20                              (merge_data_nw_2_pe[0][20]),
    .merge_valid_o_0_20                             (merge_valid_nw_2_pe[0][20]),
    .merge_ready_i_0_20                             (merge_ready_pe_2_nw[0][20]),
    .gather_data_o_0_20                             (gather_data_nw_2_pe[0][20]),
    .gather_valid_o_0_20                            (gather_valid_nw_2_pe[0][20]),
    .gather_ready_i_0_20                            (gather_ready_pe_2_nw[0][20]),
    .cast_data_i_0_21                               (cast_data_pe_2_nw[0][21]),
    .cast_valid_i_0_21                              (cast_valid_pe_2_nw[0][21]),
    .cast_ready_o_0_21                              (cast_ready_nw_2_pe[0][21]),
    .merge_data_i_0_21                              (merge_data_pe_2_nw[0][21]),
    .merge_valid_i_0_21                             (merge_valid_pe_2_nw[0][21]),
    .merge_ready_o_0_21                             (merge_ready_nw_2_pe[0][21]),
    .gather_data_i_0_21                             (gather_data_pe_2_nw[0][21]),
    .gather_valid_i_0_21                            (gather_valid_pe_2_nw[0][21]),
    .gather_ready_o_0_21                            (gather_ready_nw_2_pe[0][21]),

    .cast_data_o_0_21                               (cast_data_nw_2_pe[0][21]),
    .cast_valid_o_0_21                              (cast_valid_nw_2_pe[0][21]),
    .cast_ready_i_0_21                              (cast_ready_pe_2_nw[0][21]),
    .merge_data_o_0_21                              (merge_data_nw_2_pe[0][21]),
    .merge_valid_o_0_21                             (merge_valid_nw_2_pe[0][21]),
    .merge_ready_i_0_21                             (merge_ready_pe_2_nw[0][21]),
    .gather_data_o_0_21                             (gather_data_nw_2_pe[0][21]),
    .gather_valid_o_0_21                            (gather_valid_nw_2_pe[0][21]),
    .gather_ready_i_0_21                            (gather_ready_pe_2_nw[0][21]),
    .cast_data_i_0_22                               (cast_data_pe_2_nw[0][22]),
    .cast_valid_i_0_22                              (cast_valid_pe_2_nw[0][22]),
    .cast_ready_o_0_22                              (cast_ready_nw_2_pe[0][22]),
    .merge_data_i_0_22                              (merge_data_pe_2_nw[0][22]),
    .merge_valid_i_0_22                             (merge_valid_pe_2_nw[0][22]),
    .merge_ready_o_0_22                             (merge_ready_nw_2_pe[0][22]),
    .gather_data_i_0_22                             (gather_data_pe_2_nw[0][22]),
    .gather_valid_i_0_22                            (gather_valid_pe_2_nw[0][22]),
    .gather_ready_o_0_22                            (gather_ready_nw_2_pe[0][22]),

    .cast_data_o_0_22                               (cast_data_nw_2_pe[0][22]),
    .cast_valid_o_0_22                              (cast_valid_nw_2_pe[0][22]),
    .cast_ready_i_0_22                              (cast_ready_pe_2_nw[0][22]),
    .merge_data_o_0_22                              (merge_data_nw_2_pe[0][22]),
    .merge_valid_o_0_22                             (merge_valid_nw_2_pe[0][22]),
    .merge_ready_i_0_22                             (merge_ready_pe_2_nw[0][22]),
    .gather_data_o_0_22                             (gather_data_nw_2_pe[0][22]),
    .gather_valid_o_0_22                            (gather_valid_nw_2_pe[0][22]),
    .gather_ready_i_0_22                            (gather_ready_pe_2_nw[0][22]),
    .cast_data_i_0_23                               (cast_data_pe_2_nw[0][23]),
    .cast_valid_i_0_23                              (cast_valid_pe_2_nw[0][23]),
    .cast_ready_o_0_23                              (cast_ready_nw_2_pe[0][23]),
    .merge_data_i_0_23                              (merge_data_pe_2_nw[0][23]),
    .merge_valid_i_0_23                             (merge_valid_pe_2_nw[0][23]),
    .merge_ready_o_0_23                             (merge_ready_nw_2_pe[0][23]),
    .gather_data_i_0_23                             (gather_data_pe_2_nw[0][23]),
    .gather_valid_i_0_23                            (gather_valid_pe_2_nw[0][23]),
    .gather_ready_o_0_23                            (gather_ready_nw_2_pe[0][23]),

    .cast_data_o_0_23                               (cast_data_nw_2_pe[0][23]),
    .cast_valid_o_0_23                              (cast_valid_nw_2_pe[0][23]),
    .cast_ready_i_0_23                              (cast_ready_pe_2_nw[0][23]),
    .merge_data_o_0_23                              (merge_data_nw_2_pe[0][23]),
    .merge_valid_o_0_23                             (merge_valid_nw_2_pe[0][23]),
    .merge_ready_i_0_23                             (merge_ready_pe_2_nw[0][23]),
    .gather_data_o_0_23                             (gather_data_nw_2_pe[0][23]),
    .gather_valid_o_0_23                            (gather_valid_nw_2_pe[0][23]),
    .gather_ready_i_0_23                            (gather_ready_pe_2_nw[0][23]),
    .cast_data_i_0_24                               (cast_data_pe_2_nw[0][24]),
    .cast_valid_i_0_24                              (cast_valid_pe_2_nw[0][24]),
    .cast_ready_o_0_24                              (cast_ready_nw_2_pe[0][24]),
    .merge_data_i_0_24                              (merge_data_pe_2_nw[0][24]),
    .merge_valid_i_0_24                             (merge_valid_pe_2_nw[0][24]),
    .merge_ready_o_0_24                             (merge_ready_nw_2_pe[0][24]),
    .gather_data_i_0_24                             (gather_data_pe_2_nw[0][24]),
    .gather_valid_i_0_24                            (gather_valid_pe_2_nw[0][24]),
    .gather_ready_o_0_24                            (gather_ready_nw_2_pe[0][24]),

    .cast_data_o_0_24                               (cast_data_nw_2_pe[0][24]),
    .cast_valid_o_0_24                              (cast_valid_nw_2_pe[0][24]),
    .cast_ready_i_0_24                              (cast_ready_pe_2_nw[0][24]),
    .merge_data_o_0_24                              (merge_data_nw_2_pe[0][24]),
    .merge_valid_o_0_24                             (merge_valid_nw_2_pe[0][24]),
    .merge_ready_i_0_24                             (merge_ready_pe_2_nw[0][24]),
    .gather_data_o_0_24                             (gather_data_nw_2_pe[0][24]),
    .gather_valid_o_0_24                            (gather_valid_nw_2_pe[0][24]),
    .gather_ready_i_0_24                            (gather_ready_pe_2_nw[0][24]),
    .cast_data_i_1_0                               (cast_data_pe_2_nw[1][0]),
    .cast_valid_i_1_0                              (cast_valid_pe_2_nw[1][0]),
    .cast_ready_o_1_0                              (cast_ready_nw_2_pe[1][0]),
    .merge_data_i_1_0                              (merge_data_pe_2_nw[1][0]),
    .merge_valid_i_1_0                             (merge_valid_pe_2_nw[1][0]),
    .merge_ready_o_1_0                             (merge_ready_nw_2_pe[1][0]),
    .gather_data_i_1_0                             (gather_data_pe_2_nw[1][0]),
    .gather_valid_i_1_0                            (gather_valid_pe_2_nw[1][0]),
    .gather_ready_o_1_0                            (gather_ready_nw_2_pe[1][0]),

    .cast_data_o_1_0                               (cast_data_nw_2_pe[1][0]),
    .cast_valid_o_1_0                              (cast_valid_nw_2_pe[1][0]),
    .cast_ready_i_1_0                              (cast_ready_pe_2_nw[1][0]),
    .merge_data_o_1_0                              (merge_data_nw_2_pe[1][0]),
    .merge_valid_o_1_0                             (merge_valid_nw_2_pe[1][0]),
    .merge_ready_i_1_0                             (merge_ready_pe_2_nw[1][0]),
    .gather_data_o_1_0                             (gather_data_nw_2_pe[1][0]),
    .gather_valid_o_1_0                            (gather_valid_nw_2_pe[1][0]),
    .gather_ready_i_1_0                            (gather_ready_pe_2_nw[1][0]),
    .cast_data_i_1_1                               (cast_data_pe_2_nw[1][1]),
    .cast_valid_i_1_1                              (cast_valid_pe_2_nw[1][1]),
    .cast_ready_o_1_1                              (cast_ready_nw_2_pe[1][1]),
    .merge_data_i_1_1                              (merge_data_pe_2_nw[1][1]),
    .merge_valid_i_1_1                             (merge_valid_pe_2_nw[1][1]),
    .merge_ready_o_1_1                             (merge_ready_nw_2_pe[1][1]),
    .gather_data_i_1_1                             (gather_data_pe_2_nw[1][1]),
    .gather_valid_i_1_1                            (gather_valid_pe_2_nw[1][1]),
    .gather_ready_o_1_1                            (gather_ready_nw_2_pe[1][1]),

    .cast_data_o_1_1                               (cast_data_nw_2_pe[1][1]),
    .cast_valid_o_1_1                              (cast_valid_nw_2_pe[1][1]),
    .cast_ready_i_1_1                              (cast_ready_pe_2_nw[1][1]),
    .merge_data_o_1_1                              (merge_data_nw_2_pe[1][1]),
    .merge_valid_o_1_1                             (merge_valid_nw_2_pe[1][1]),
    .merge_ready_i_1_1                             (merge_ready_pe_2_nw[1][1]),
    .gather_data_o_1_1                             (gather_data_nw_2_pe[1][1]),
    .gather_valid_o_1_1                            (gather_valid_nw_2_pe[1][1]),
    .gather_ready_i_1_1                            (gather_ready_pe_2_nw[1][1]),
    .cast_data_i_1_2                               (cast_data_pe_2_nw[1][2]),
    .cast_valid_i_1_2                              (cast_valid_pe_2_nw[1][2]),
    .cast_ready_o_1_2                              (cast_ready_nw_2_pe[1][2]),
    .merge_data_i_1_2                              (merge_data_pe_2_nw[1][2]),
    .merge_valid_i_1_2                             (merge_valid_pe_2_nw[1][2]),
    .merge_ready_o_1_2                             (merge_ready_nw_2_pe[1][2]),
    .gather_data_i_1_2                             (gather_data_pe_2_nw[1][2]),
    .gather_valid_i_1_2                            (gather_valid_pe_2_nw[1][2]),
    .gather_ready_o_1_2                            (gather_ready_nw_2_pe[1][2]),

    .cast_data_o_1_2                               (cast_data_nw_2_pe[1][2]),
    .cast_valid_o_1_2                              (cast_valid_nw_2_pe[1][2]),
    .cast_ready_i_1_2                              (cast_ready_pe_2_nw[1][2]),
    .merge_data_o_1_2                              (merge_data_nw_2_pe[1][2]),
    .merge_valid_o_1_2                             (merge_valid_nw_2_pe[1][2]),
    .merge_ready_i_1_2                             (merge_ready_pe_2_nw[1][2]),
    .gather_data_o_1_2                             (gather_data_nw_2_pe[1][2]),
    .gather_valid_o_1_2                            (gather_valid_nw_2_pe[1][2]),
    .gather_ready_i_1_2                            (gather_ready_pe_2_nw[1][2]),
    .cast_data_i_1_3                               (cast_data_pe_2_nw[1][3]),
    .cast_valid_i_1_3                              (cast_valid_pe_2_nw[1][3]),
    .cast_ready_o_1_3                              (cast_ready_nw_2_pe[1][3]),
    .merge_data_i_1_3                              (merge_data_pe_2_nw[1][3]),
    .merge_valid_i_1_3                             (merge_valid_pe_2_nw[1][3]),
    .merge_ready_o_1_3                             (merge_ready_nw_2_pe[1][3]),
    .gather_data_i_1_3                             (gather_data_pe_2_nw[1][3]),
    .gather_valid_i_1_3                            (gather_valid_pe_2_nw[1][3]),
    .gather_ready_o_1_3                            (gather_ready_nw_2_pe[1][3]),

    .cast_data_o_1_3                               (cast_data_nw_2_pe[1][3]),
    .cast_valid_o_1_3                              (cast_valid_nw_2_pe[1][3]),
    .cast_ready_i_1_3                              (cast_ready_pe_2_nw[1][3]),
    .merge_data_o_1_3                              (merge_data_nw_2_pe[1][3]),
    .merge_valid_o_1_3                             (merge_valid_nw_2_pe[1][3]),
    .merge_ready_i_1_3                             (merge_ready_pe_2_nw[1][3]),
    .gather_data_o_1_3                             (gather_data_nw_2_pe[1][3]),
    .gather_valid_o_1_3                            (gather_valid_nw_2_pe[1][3]),
    .gather_ready_i_1_3                            (gather_ready_pe_2_nw[1][3]),
    .cast_data_i_1_4                               (cast_data_pe_2_nw[1][4]),
    .cast_valid_i_1_4                              (cast_valid_pe_2_nw[1][4]),
    .cast_ready_o_1_4                              (cast_ready_nw_2_pe[1][4]),
    .merge_data_i_1_4                              (merge_data_pe_2_nw[1][4]),
    .merge_valid_i_1_4                             (merge_valid_pe_2_nw[1][4]),
    .merge_ready_o_1_4                             (merge_ready_nw_2_pe[1][4]),
    .gather_data_i_1_4                             (gather_data_pe_2_nw[1][4]),
    .gather_valid_i_1_4                            (gather_valid_pe_2_nw[1][4]),
    .gather_ready_o_1_4                            (gather_ready_nw_2_pe[1][4]),

    .cast_data_o_1_4                               (cast_data_nw_2_pe[1][4]),
    .cast_valid_o_1_4                              (cast_valid_nw_2_pe[1][4]),
    .cast_ready_i_1_4                              (cast_ready_pe_2_nw[1][4]),
    .merge_data_o_1_4                              (merge_data_nw_2_pe[1][4]),
    .merge_valid_o_1_4                             (merge_valid_nw_2_pe[1][4]),
    .merge_ready_i_1_4                             (merge_ready_pe_2_nw[1][4]),
    .gather_data_o_1_4                             (gather_data_nw_2_pe[1][4]),
    .gather_valid_o_1_4                            (gather_valid_nw_2_pe[1][4]),
    .gather_ready_i_1_4                            (gather_ready_pe_2_nw[1][4]),
    .cast_data_i_1_5                               (cast_data_pe_2_nw[1][5]),
    .cast_valid_i_1_5                              (cast_valid_pe_2_nw[1][5]),
    .cast_ready_o_1_5                              (cast_ready_nw_2_pe[1][5]),
    .merge_data_i_1_5                              (merge_data_pe_2_nw[1][5]),
    .merge_valid_i_1_5                             (merge_valid_pe_2_nw[1][5]),
    .merge_ready_o_1_5                             (merge_ready_nw_2_pe[1][5]),
    .gather_data_i_1_5                             (gather_data_pe_2_nw[1][5]),
    .gather_valid_i_1_5                            (gather_valid_pe_2_nw[1][5]),
    .gather_ready_o_1_5                            (gather_ready_nw_2_pe[1][5]),

    .cast_data_o_1_5                               (cast_data_nw_2_pe[1][5]),
    .cast_valid_o_1_5                              (cast_valid_nw_2_pe[1][5]),
    .cast_ready_i_1_5                              (cast_ready_pe_2_nw[1][5]),
    .merge_data_o_1_5                              (merge_data_nw_2_pe[1][5]),
    .merge_valid_o_1_5                             (merge_valid_nw_2_pe[1][5]),
    .merge_ready_i_1_5                             (merge_ready_pe_2_nw[1][5]),
    .gather_data_o_1_5                             (gather_data_nw_2_pe[1][5]),
    .gather_valid_o_1_5                            (gather_valid_nw_2_pe[1][5]),
    .gather_ready_i_1_5                            (gather_ready_pe_2_nw[1][5]),
    .cast_data_i_1_6                               (cast_data_pe_2_nw[1][6]),
    .cast_valid_i_1_6                              (cast_valid_pe_2_nw[1][6]),
    .cast_ready_o_1_6                              (cast_ready_nw_2_pe[1][6]),
    .merge_data_i_1_6                              (merge_data_pe_2_nw[1][6]),
    .merge_valid_i_1_6                             (merge_valid_pe_2_nw[1][6]),
    .merge_ready_o_1_6                             (merge_ready_nw_2_pe[1][6]),
    .gather_data_i_1_6                             (gather_data_pe_2_nw[1][6]),
    .gather_valid_i_1_6                            (gather_valid_pe_2_nw[1][6]),
    .gather_ready_o_1_6                            (gather_ready_nw_2_pe[1][6]),

    .cast_data_o_1_6                               (cast_data_nw_2_pe[1][6]),
    .cast_valid_o_1_6                              (cast_valid_nw_2_pe[1][6]),
    .cast_ready_i_1_6                              (cast_ready_pe_2_nw[1][6]),
    .merge_data_o_1_6                              (merge_data_nw_2_pe[1][6]),
    .merge_valid_o_1_6                             (merge_valid_nw_2_pe[1][6]),
    .merge_ready_i_1_6                             (merge_ready_pe_2_nw[1][6]),
    .gather_data_o_1_6                             (gather_data_nw_2_pe[1][6]),
    .gather_valid_o_1_6                            (gather_valid_nw_2_pe[1][6]),
    .gather_ready_i_1_6                            (gather_ready_pe_2_nw[1][6]),
    .cast_data_i_1_7                               (cast_data_pe_2_nw[1][7]),
    .cast_valid_i_1_7                              (cast_valid_pe_2_nw[1][7]),
    .cast_ready_o_1_7                              (cast_ready_nw_2_pe[1][7]),
    .merge_data_i_1_7                              (merge_data_pe_2_nw[1][7]),
    .merge_valid_i_1_7                             (merge_valid_pe_2_nw[1][7]),
    .merge_ready_o_1_7                             (merge_ready_nw_2_pe[1][7]),
    .gather_data_i_1_7                             (gather_data_pe_2_nw[1][7]),
    .gather_valid_i_1_7                            (gather_valid_pe_2_nw[1][7]),
    .gather_ready_o_1_7                            (gather_ready_nw_2_pe[1][7]),

    .cast_data_o_1_7                               (cast_data_nw_2_pe[1][7]),
    .cast_valid_o_1_7                              (cast_valid_nw_2_pe[1][7]),
    .cast_ready_i_1_7                              (cast_ready_pe_2_nw[1][7]),
    .merge_data_o_1_7                              (merge_data_nw_2_pe[1][7]),
    .merge_valid_o_1_7                             (merge_valid_nw_2_pe[1][7]),
    .merge_ready_i_1_7                             (merge_ready_pe_2_nw[1][7]),
    .gather_data_o_1_7                             (gather_data_nw_2_pe[1][7]),
    .gather_valid_o_1_7                            (gather_valid_nw_2_pe[1][7]),
    .gather_ready_i_1_7                            (gather_ready_pe_2_nw[1][7]),
    .cast_data_i_1_8                               (cast_data_pe_2_nw[1][8]),
    .cast_valid_i_1_8                              (cast_valid_pe_2_nw[1][8]),
    .cast_ready_o_1_8                              (cast_ready_nw_2_pe[1][8]),
    .merge_data_i_1_8                              (merge_data_pe_2_nw[1][8]),
    .merge_valid_i_1_8                             (merge_valid_pe_2_nw[1][8]),
    .merge_ready_o_1_8                             (merge_ready_nw_2_pe[1][8]),
    .gather_data_i_1_8                             (gather_data_pe_2_nw[1][8]),
    .gather_valid_i_1_8                            (gather_valid_pe_2_nw[1][8]),
    .gather_ready_o_1_8                            (gather_ready_nw_2_pe[1][8]),

    .cast_data_o_1_8                               (cast_data_nw_2_pe[1][8]),
    .cast_valid_o_1_8                              (cast_valid_nw_2_pe[1][8]),
    .cast_ready_i_1_8                              (cast_ready_pe_2_nw[1][8]),
    .merge_data_o_1_8                              (merge_data_nw_2_pe[1][8]),
    .merge_valid_o_1_8                             (merge_valid_nw_2_pe[1][8]),
    .merge_ready_i_1_8                             (merge_ready_pe_2_nw[1][8]),
    .gather_data_o_1_8                             (gather_data_nw_2_pe[1][8]),
    .gather_valid_o_1_8                            (gather_valid_nw_2_pe[1][8]),
    .gather_ready_i_1_8                            (gather_ready_pe_2_nw[1][8]),
    .cast_data_i_1_9                               (cast_data_pe_2_nw[1][9]),
    .cast_valid_i_1_9                              (cast_valid_pe_2_nw[1][9]),
    .cast_ready_o_1_9                              (cast_ready_nw_2_pe[1][9]),
    .merge_data_i_1_9                              (merge_data_pe_2_nw[1][9]),
    .merge_valid_i_1_9                             (merge_valid_pe_2_nw[1][9]),
    .merge_ready_o_1_9                             (merge_ready_nw_2_pe[1][9]),
    .gather_data_i_1_9                             (gather_data_pe_2_nw[1][9]),
    .gather_valid_i_1_9                            (gather_valid_pe_2_nw[1][9]),
    .gather_ready_o_1_9                            (gather_ready_nw_2_pe[1][9]),

    .cast_data_o_1_9                               (cast_data_nw_2_pe[1][9]),
    .cast_valid_o_1_9                              (cast_valid_nw_2_pe[1][9]),
    .cast_ready_i_1_9                              (cast_ready_pe_2_nw[1][9]),
    .merge_data_o_1_9                              (merge_data_nw_2_pe[1][9]),
    .merge_valid_o_1_9                             (merge_valid_nw_2_pe[1][9]),
    .merge_ready_i_1_9                             (merge_ready_pe_2_nw[1][9]),
    .gather_data_o_1_9                             (gather_data_nw_2_pe[1][9]),
    .gather_valid_o_1_9                            (gather_valid_nw_2_pe[1][9]),
    .gather_ready_i_1_9                            (gather_ready_pe_2_nw[1][9]),
    .cast_data_i_1_10                               (cast_data_pe_2_nw[1][10]),
    .cast_valid_i_1_10                              (cast_valid_pe_2_nw[1][10]),
    .cast_ready_o_1_10                              (cast_ready_nw_2_pe[1][10]),
    .merge_data_i_1_10                              (merge_data_pe_2_nw[1][10]),
    .merge_valid_i_1_10                             (merge_valid_pe_2_nw[1][10]),
    .merge_ready_o_1_10                             (merge_ready_nw_2_pe[1][10]),
    .gather_data_i_1_10                             (gather_data_pe_2_nw[1][10]),
    .gather_valid_i_1_10                            (gather_valid_pe_2_nw[1][10]),
    .gather_ready_o_1_10                            (gather_ready_nw_2_pe[1][10]),

    .cast_data_o_1_10                               (cast_data_nw_2_pe[1][10]),
    .cast_valid_o_1_10                              (cast_valid_nw_2_pe[1][10]),
    .cast_ready_i_1_10                              (cast_ready_pe_2_nw[1][10]),
    .merge_data_o_1_10                              (merge_data_nw_2_pe[1][10]),
    .merge_valid_o_1_10                             (merge_valid_nw_2_pe[1][10]),
    .merge_ready_i_1_10                             (merge_ready_pe_2_nw[1][10]),
    .gather_data_o_1_10                             (gather_data_nw_2_pe[1][10]),
    .gather_valid_o_1_10                            (gather_valid_nw_2_pe[1][10]),
    .gather_ready_i_1_10                            (gather_ready_pe_2_nw[1][10]),
    .cast_data_i_1_11                               (cast_data_pe_2_nw[1][11]),
    .cast_valid_i_1_11                              (cast_valid_pe_2_nw[1][11]),
    .cast_ready_o_1_11                              (cast_ready_nw_2_pe[1][11]),
    .merge_data_i_1_11                              (merge_data_pe_2_nw[1][11]),
    .merge_valid_i_1_11                             (merge_valid_pe_2_nw[1][11]),
    .merge_ready_o_1_11                             (merge_ready_nw_2_pe[1][11]),
    .gather_data_i_1_11                             (gather_data_pe_2_nw[1][11]),
    .gather_valid_i_1_11                            (gather_valid_pe_2_nw[1][11]),
    .gather_ready_o_1_11                            (gather_ready_nw_2_pe[1][11]),

    .cast_data_o_1_11                               (cast_data_nw_2_pe[1][11]),
    .cast_valid_o_1_11                              (cast_valid_nw_2_pe[1][11]),
    .cast_ready_i_1_11                              (cast_ready_pe_2_nw[1][11]),
    .merge_data_o_1_11                              (merge_data_nw_2_pe[1][11]),
    .merge_valid_o_1_11                             (merge_valid_nw_2_pe[1][11]),
    .merge_ready_i_1_11                             (merge_ready_pe_2_nw[1][11]),
    .gather_data_o_1_11                             (gather_data_nw_2_pe[1][11]),
    .gather_valid_o_1_11                            (gather_valid_nw_2_pe[1][11]),
    .gather_ready_i_1_11                            (gather_ready_pe_2_nw[1][11]),
    .cast_data_i_1_12                               (cast_data_pe_2_nw[1][12]),
    .cast_valid_i_1_12                              (cast_valid_pe_2_nw[1][12]),
    .cast_ready_o_1_12                              (cast_ready_nw_2_pe[1][12]),
    .merge_data_i_1_12                              (merge_data_pe_2_nw[1][12]),
    .merge_valid_i_1_12                             (merge_valid_pe_2_nw[1][12]),
    .merge_ready_o_1_12                             (merge_ready_nw_2_pe[1][12]),
    .gather_data_i_1_12                             (gather_data_pe_2_nw[1][12]),
    .gather_valid_i_1_12                            (gather_valid_pe_2_nw[1][12]),
    .gather_ready_o_1_12                            (gather_ready_nw_2_pe[1][12]),

    .cast_data_o_1_12                               (cast_data_nw_2_pe[1][12]),
    .cast_valid_o_1_12                              (cast_valid_nw_2_pe[1][12]),
    .cast_ready_i_1_12                              (cast_ready_pe_2_nw[1][12]),
    .merge_data_o_1_12                              (merge_data_nw_2_pe[1][12]),
    .merge_valid_o_1_12                             (merge_valid_nw_2_pe[1][12]),
    .merge_ready_i_1_12                             (merge_ready_pe_2_nw[1][12]),
    .gather_data_o_1_12                             (gather_data_nw_2_pe[1][12]),
    .gather_valid_o_1_12                            (gather_valid_nw_2_pe[1][12]),
    .gather_ready_i_1_12                            (gather_ready_pe_2_nw[1][12]),
    .cast_data_i_1_13                               (cast_data_pe_2_nw[1][13]),
    .cast_valid_i_1_13                              (cast_valid_pe_2_nw[1][13]),
    .cast_ready_o_1_13                              (cast_ready_nw_2_pe[1][13]),
    .merge_data_i_1_13                              (merge_data_pe_2_nw[1][13]),
    .merge_valid_i_1_13                             (merge_valid_pe_2_nw[1][13]),
    .merge_ready_o_1_13                             (merge_ready_nw_2_pe[1][13]),
    .gather_data_i_1_13                             (gather_data_pe_2_nw[1][13]),
    .gather_valid_i_1_13                            (gather_valid_pe_2_nw[1][13]),
    .gather_ready_o_1_13                            (gather_ready_nw_2_pe[1][13]),

    .cast_data_o_1_13                               (cast_data_nw_2_pe[1][13]),
    .cast_valid_o_1_13                              (cast_valid_nw_2_pe[1][13]),
    .cast_ready_i_1_13                              (cast_ready_pe_2_nw[1][13]),
    .merge_data_o_1_13                              (merge_data_nw_2_pe[1][13]),
    .merge_valid_o_1_13                             (merge_valid_nw_2_pe[1][13]),
    .merge_ready_i_1_13                             (merge_ready_pe_2_nw[1][13]),
    .gather_data_o_1_13                             (gather_data_nw_2_pe[1][13]),
    .gather_valid_o_1_13                            (gather_valid_nw_2_pe[1][13]),
    .gather_ready_i_1_13                            (gather_ready_pe_2_nw[1][13]),
    .cast_data_i_1_14                               (cast_data_pe_2_nw[1][14]),
    .cast_valid_i_1_14                              (cast_valid_pe_2_nw[1][14]),
    .cast_ready_o_1_14                              (cast_ready_nw_2_pe[1][14]),
    .merge_data_i_1_14                              (merge_data_pe_2_nw[1][14]),
    .merge_valid_i_1_14                             (merge_valid_pe_2_nw[1][14]),
    .merge_ready_o_1_14                             (merge_ready_nw_2_pe[1][14]),
    .gather_data_i_1_14                             (gather_data_pe_2_nw[1][14]),
    .gather_valid_i_1_14                            (gather_valid_pe_2_nw[1][14]),
    .gather_ready_o_1_14                            (gather_ready_nw_2_pe[1][14]),

    .cast_data_o_1_14                               (cast_data_nw_2_pe[1][14]),
    .cast_valid_o_1_14                              (cast_valid_nw_2_pe[1][14]),
    .cast_ready_i_1_14                              (cast_ready_pe_2_nw[1][14]),
    .merge_data_o_1_14                              (merge_data_nw_2_pe[1][14]),
    .merge_valid_o_1_14                             (merge_valid_nw_2_pe[1][14]),
    .merge_ready_i_1_14                             (merge_ready_pe_2_nw[1][14]),
    .gather_data_o_1_14                             (gather_data_nw_2_pe[1][14]),
    .gather_valid_o_1_14                            (gather_valid_nw_2_pe[1][14]),
    .gather_ready_i_1_14                            (gather_ready_pe_2_nw[1][14]),
    .cast_data_i_1_15                               (cast_data_pe_2_nw[1][15]),
    .cast_valid_i_1_15                              (cast_valid_pe_2_nw[1][15]),
    .cast_ready_o_1_15                              (cast_ready_nw_2_pe[1][15]),
    .merge_data_i_1_15                              (merge_data_pe_2_nw[1][15]),
    .merge_valid_i_1_15                             (merge_valid_pe_2_nw[1][15]),
    .merge_ready_o_1_15                             (merge_ready_nw_2_pe[1][15]),
    .gather_data_i_1_15                             (gather_data_pe_2_nw[1][15]),
    .gather_valid_i_1_15                            (gather_valid_pe_2_nw[1][15]),
    .gather_ready_o_1_15                            (gather_ready_nw_2_pe[1][15]),

    .cast_data_o_1_15                               (cast_data_nw_2_pe[1][15]),
    .cast_valid_o_1_15                              (cast_valid_nw_2_pe[1][15]),
    .cast_ready_i_1_15                              (cast_ready_pe_2_nw[1][15]),
    .merge_data_o_1_15                              (merge_data_nw_2_pe[1][15]),
    .merge_valid_o_1_15                             (merge_valid_nw_2_pe[1][15]),
    .merge_ready_i_1_15                             (merge_ready_pe_2_nw[1][15]),
    .gather_data_o_1_15                             (gather_data_nw_2_pe[1][15]),
    .gather_valid_o_1_15                            (gather_valid_nw_2_pe[1][15]),
    .gather_ready_i_1_15                            (gather_ready_pe_2_nw[1][15]),
    .cast_data_i_1_16                               (cast_data_pe_2_nw[1][16]),
    .cast_valid_i_1_16                              (cast_valid_pe_2_nw[1][16]),
    .cast_ready_o_1_16                              (cast_ready_nw_2_pe[1][16]),
    .merge_data_i_1_16                              (merge_data_pe_2_nw[1][16]),
    .merge_valid_i_1_16                             (merge_valid_pe_2_nw[1][16]),
    .merge_ready_o_1_16                             (merge_ready_nw_2_pe[1][16]),
    .gather_data_i_1_16                             (gather_data_pe_2_nw[1][16]),
    .gather_valid_i_1_16                            (gather_valid_pe_2_nw[1][16]),
    .gather_ready_o_1_16                            (gather_ready_nw_2_pe[1][16]),

    .cast_data_o_1_16                               (cast_data_nw_2_pe[1][16]),
    .cast_valid_o_1_16                              (cast_valid_nw_2_pe[1][16]),
    .cast_ready_i_1_16                              (cast_ready_pe_2_nw[1][16]),
    .merge_data_o_1_16                              (merge_data_nw_2_pe[1][16]),
    .merge_valid_o_1_16                             (merge_valid_nw_2_pe[1][16]),
    .merge_ready_i_1_16                             (merge_ready_pe_2_nw[1][16]),
    .gather_data_o_1_16                             (gather_data_nw_2_pe[1][16]),
    .gather_valid_o_1_16                            (gather_valid_nw_2_pe[1][16]),
    .gather_ready_i_1_16                            (gather_ready_pe_2_nw[1][16]),
    .cast_data_i_1_17                               (cast_data_pe_2_nw[1][17]),
    .cast_valid_i_1_17                              (cast_valid_pe_2_nw[1][17]),
    .cast_ready_o_1_17                              (cast_ready_nw_2_pe[1][17]),
    .merge_data_i_1_17                              (merge_data_pe_2_nw[1][17]),
    .merge_valid_i_1_17                             (merge_valid_pe_2_nw[1][17]),
    .merge_ready_o_1_17                             (merge_ready_nw_2_pe[1][17]),
    .gather_data_i_1_17                             (gather_data_pe_2_nw[1][17]),
    .gather_valid_i_1_17                            (gather_valid_pe_2_nw[1][17]),
    .gather_ready_o_1_17                            (gather_ready_nw_2_pe[1][17]),

    .cast_data_o_1_17                               (cast_data_nw_2_pe[1][17]),
    .cast_valid_o_1_17                              (cast_valid_nw_2_pe[1][17]),
    .cast_ready_i_1_17                              (cast_ready_pe_2_nw[1][17]),
    .merge_data_o_1_17                              (merge_data_nw_2_pe[1][17]),
    .merge_valid_o_1_17                             (merge_valid_nw_2_pe[1][17]),
    .merge_ready_i_1_17                             (merge_ready_pe_2_nw[1][17]),
    .gather_data_o_1_17                             (gather_data_nw_2_pe[1][17]),
    .gather_valid_o_1_17                            (gather_valid_nw_2_pe[1][17]),
    .gather_ready_i_1_17                            (gather_ready_pe_2_nw[1][17]),
    .cast_data_i_1_18                               (cast_data_pe_2_nw[1][18]),
    .cast_valid_i_1_18                              (cast_valid_pe_2_nw[1][18]),
    .cast_ready_o_1_18                              (cast_ready_nw_2_pe[1][18]),
    .merge_data_i_1_18                              (merge_data_pe_2_nw[1][18]),
    .merge_valid_i_1_18                             (merge_valid_pe_2_nw[1][18]),
    .merge_ready_o_1_18                             (merge_ready_nw_2_pe[1][18]),
    .gather_data_i_1_18                             (gather_data_pe_2_nw[1][18]),
    .gather_valid_i_1_18                            (gather_valid_pe_2_nw[1][18]),
    .gather_ready_o_1_18                            (gather_ready_nw_2_pe[1][18]),

    .cast_data_o_1_18                               (cast_data_nw_2_pe[1][18]),
    .cast_valid_o_1_18                              (cast_valid_nw_2_pe[1][18]),
    .cast_ready_i_1_18                              (cast_ready_pe_2_nw[1][18]),
    .merge_data_o_1_18                              (merge_data_nw_2_pe[1][18]),
    .merge_valid_o_1_18                             (merge_valid_nw_2_pe[1][18]),
    .merge_ready_i_1_18                             (merge_ready_pe_2_nw[1][18]),
    .gather_data_o_1_18                             (gather_data_nw_2_pe[1][18]),
    .gather_valid_o_1_18                            (gather_valid_nw_2_pe[1][18]),
    .gather_ready_i_1_18                            (gather_ready_pe_2_nw[1][18]),
    .cast_data_i_1_19                               (cast_data_pe_2_nw[1][19]),
    .cast_valid_i_1_19                              (cast_valid_pe_2_nw[1][19]),
    .cast_ready_o_1_19                              (cast_ready_nw_2_pe[1][19]),
    .merge_data_i_1_19                              (merge_data_pe_2_nw[1][19]),
    .merge_valid_i_1_19                             (merge_valid_pe_2_nw[1][19]),
    .merge_ready_o_1_19                             (merge_ready_nw_2_pe[1][19]),
    .gather_data_i_1_19                             (gather_data_pe_2_nw[1][19]),
    .gather_valid_i_1_19                            (gather_valid_pe_2_nw[1][19]),
    .gather_ready_o_1_19                            (gather_ready_nw_2_pe[1][19]),

    .cast_data_o_1_19                               (cast_data_nw_2_pe[1][19]),
    .cast_valid_o_1_19                              (cast_valid_nw_2_pe[1][19]),
    .cast_ready_i_1_19                              (cast_ready_pe_2_nw[1][19]),
    .merge_data_o_1_19                              (merge_data_nw_2_pe[1][19]),
    .merge_valid_o_1_19                             (merge_valid_nw_2_pe[1][19]),
    .merge_ready_i_1_19                             (merge_ready_pe_2_nw[1][19]),
    .gather_data_o_1_19                             (gather_data_nw_2_pe[1][19]),
    .gather_valid_o_1_19                            (gather_valid_nw_2_pe[1][19]),
    .gather_ready_i_1_19                            (gather_ready_pe_2_nw[1][19]),
    .cast_data_i_1_20                               (cast_data_pe_2_nw[1][20]),
    .cast_valid_i_1_20                              (cast_valid_pe_2_nw[1][20]),
    .cast_ready_o_1_20                              (cast_ready_nw_2_pe[1][20]),
    .merge_data_i_1_20                              (merge_data_pe_2_nw[1][20]),
    .merge_valid_i_1_20                             (merge_valid_pe_2_nw[1][20]),
    .merge_ready_o_1_20                             (merge_ready_nw_2_pe[1][20]),
    .gather_data_i_1_20                             (gather_data_pe_2_nw[1][20]),
    .gather_valid_i_1_20                            (gather_valid_pe_2_nw[1][20]),
    .gather_ready_o_1_20                            (gather_ready_nw_2_pe[1][20]),

    .cast_data_o_1_20                               (cast_data_nw_2_pe[1][20]),
    .cast_valid_o_1_20                              (cast_valid_nw_2_pe[1][20]),
    .cast_ready_i_1_20                              (cast_ready_pe_2_nw[1][20]),
    .merge_data_o_1_20                              (merge_data_nw_2_pe[1][20]),
    .merge_valid_o_1_20                             (merge_valid_nw_2_pe[1][20]),
    .merge_ready_i_1_20                             (merge_ready_pe_2_nw[1][20]),
    .gather_data_o_1_20                             (gather_data_nw_2_pe[1][20]),
    .gather_valid_o_1_20                            (gather_valid_nw_2_pe[1][20]),
    .gather_ready_i_1_20                            (gather_ready_pe_2_nw[1][20]),
    .cast_data_i_1_21                               (cast_data_pe_2_nw[1][21]),
    .cast_valid_i_1_21                              (cast_valid_pe_2_nw[1][21]),
    .cast_ready_o_1_21                              (cast_ready_nw_2_pe[1][21]),
    .merge_data_i_1_21                              (merge_data_pe_2_nw[1][21]),
    .merge_valid_i_1_21                             (merge_valid_pe_2_nw[1][21]),
    .merge_ready_o_1_21                             (merge_ready_nw_2_pe[1][21]),
    .gather_data_i_1_21                             (gather_data_pe_2_nw[1][21]),
    .gather_valid_i_1_21                            (gather_valid_pe_2_nw[1][21]),
    .gather_ready_o_1_21                            (gather_ready_nw_2_pe[1][21]),

    .cast_data_o_1_21                               (cast_data_nw_2_pe[1][21]),
    .cast_valid_o_1_21                              (cast_valid_nw_2_pe[1][21]),
    .cast_ready_i_1_21                              (cast_ready_pe_2_nw[1][21]),
    .merge_data_o_1_21                              (merge_data_nw_2_pe[1][21]),
    .merge_valid_o_1_21                             (merge_valid_nw_2_pe[1][21]),
    .merge_ready_i_1_21                             (merge_ready_pe_2_nw[1][21]),
    .gather_data_o_1_21                             (gather_data_nw_2_pe[1][21]),
    .gather_valid_o_1_21                            (gather_valid_nw_2_pe[1][21]),
    .gather_ready_i_1_21                            (gather_ready_pe_2_nw[1][21]),
    .cast_data_i_1_22                               (cast_data_pe_2_nw[1][22]),
    .cast_valid_i_1_22                              (cast_valid_pe_2_nw[1][22]),
    .cast_ready_o_1_22                              (cast_ready_nw_2_pe[1][22]),
    .merge_data_i_1_22                              (merge_data_pe_2_nw[1][22]),
    .merge_valid_i_1_22                             (merge_valid_pe_2_nw[1][22]),
    .merge_ready_o_1_22                             (merge_ready_nw_2_pe[1][22]),
    .gather_data_i_1_22                             (gather_data_pe_2_nw[1][22]),
    .gather_valid_i_1_22                            (gather_valid_pe_2_nw[1][22]),
    .gather_ready_o_1_22                            (gather_ready_nw_2_pe[1][22]),

    .cast_data_o_1_22                               (cast_data_nw_2_pe[1][22]),
    .cast_valid_o_1_22                              (cast_valid_nw_2_pe[1][22]),
    .cast_ready_i_1_22                              (cast_ready_pe_2_nw[1][22]),
    .merge_data_o_1_22                              (merge_data_nw_2_pe[1][22]),
    .merge_valid_o_1_22                             (merge_valid_nw_2_pe[1][22]),
    .merge_ready_i_1_22                             (merge_ready_pe_2_nw[1][22]),
    .gather_data_o_1_22                             (gather_data_nw_2_pe[1][22]),
    .gather_valid_o_1_22                            (gather_valid_nw_2_pe[1][22]),
    .gather_ready_i_1_22                            (gather_ready_pe_2_nw[1][22]),
    .cast_data_i_1_23                               (cast_data_pe_2_nw[1][23]),
    .cast_valid_i_1_23                              (cast_valid_pe_2_nw[1][23]),
    .cast_ready_o_1_23                              (cast_ready_nw_2_pe[1][23]),
    .merge_data_i_1_23                              (merge_data_pe_2_nw[1][23]),
    .merge_valid_i_1_23                             (merge_valid_pe_2_nw[1][23]),
    .merge_ready_o_1_23                             (merge_ready_nw_2_pe[1][23]),
    .gather_data_i_1_23                             (gather_data_pe_2_nw[1][23]),
    .gather_valid_i_1_23                            (gather_valid_pe_2_nw[1][23]),
    .gather_ready_o_1_23                            (gather_ready_nw_2_pe[1][23]),

    .cast_data_o_1_23                               (cast_data_nw_2_pe[1][23]),
    .cast_valid_o_1_23                              (cast_valid_nw_2_pe[1][23]),
    .cast_ready_i_1_23                              (cast_ready_pe_2_nw[1][23]),
    .merge_data_o_1_23                              (merge_data_nw_2_pe[1][23]),
    .merge_valid_o_1_23                             (merge_valid_nw_2_pe[1][23]),
    .merge_ready_i_1_23                             (merge_ready_pe_2_nw[1][23]),
    .gather_data_o_1_23                             (gather_data_nw_2_pe[1][23]),
    .gather_valid_o_1_23                            (gather_valid_nw_2_pe[1][23]),
    .gather_ready_i_1_23                            (gather_ready_pe_2_nw[1][23]),
    .cast_data_i_1_24                               (cast_data_pe_2_nw[1][24]),
    .cast_valid_i_1_24                              (cast_valid_pe_2_nw[1][24]),
    .cast_ready_o_1_24                              (cast_ready_nw_2_pe[1][24]),
    .merge_data_i_1_24                              (merge_data_pe_2_nw[1][24]),
    .merge_valid_i_1_24                             (merge_valid_pe_2_nw[1][24]),
    .merge_ready_o_1_24                             (merge_ready_nw_2_pe[1][24]),
    .gather_data_i_1_24                             (gather_data_pe_2_nw[1][24]),
    .gather_valid_i_1_24                            (gather_valid_pe_2_nw[1][24]),
    .gather_ready_o_1_24                            (gather_ready_nw_2_pe[1][24]),

    .cast_data_o_1_24                               (cast_data_nw_2_pe[1][24]),
    .cast_valid_o_1_24                              (cast_valid_nw_2_pe[1][24]),
    .cast_ready_i_1_24                              (cast_ready_pe_2_nw[1][24]),
    .merge_data_o_1_24                              (merge_data_nw_2_pe[1][24]),
    .merge_valid_o_1_24                             (merge_valid_nw_2_pe[1][24]),
    .merge_ready_i_1_24                             (merge_ready_pe_2_nw[1][24]),
    .gather_data_o_1_24                             (gather_data_nw_2_pe[1][24]),
    .gather_valid_o_1_24                            (gather_valid_nw_2_pe[1][24]),
    .gather_ready_i_1_24                            (gather_ready_pe_2_nw[1][24]),
    .cast_data_i_2_0                               (cast_data_pe_2_nw[2][0]),
    .cast_valid_i_2_0                              (cast_valid_pe_2_nw[2][0]),
    .cast_ready_o_2_0                              (cast_ready_nw_2_pe[2][0]),
    .merge_data_i_2_0                              (merge_data_pe_2_nw[2][0]),
    .merge_valid_i_2_0                             (merge_valid_pe_2_nw[2][0]),
    .merge_ready_o_2_0                             (merge_ready_nw_2_pe[2][0]),
    .gather_data_i_2_0                             (gather_data_pe_2_nw[2][0]),
    .gather_valid_i_2_0                            (gather_valid_pe_2_nw[2][0]),
    .gather_ready_o_2_0                            (gather_ready_nw_2_pe[2][0]),

    .cast_data_o_2_0                               (cast_data_nw_2_pe[2][0]),
    .cast_valid_o_2_0                              (cast_valid_nw_2_pe[2][0]),
    .cast_ready_i_2_0                              (cast_ready_pe_2_nw[2][0]),
    .merge_data_o_2_0                              (merge_data_nw_2_pe[2][0]),
    .merge_valid_o_2_0                             (merge_valid_nw_2_pe[2][0]),
    .merge_ready_i_2_0                             (merge_ready_pe_2_nw[2][0]),
    .gather_data_o_2_0                             (gather_data_nw_2_pe[2][0]),
    .gather_valid_o_2_0                            (gather_valid_nw_2_pe[2][0]),
    .gather_ready_i_2_0                            (gather_ready_pe_2_nw[2][0]),
    .cast_data_i_2_1                               (cast_data_pe_2_nw[2][1]),
    .cast_valid_i_2_1                              (cast_valid_pe_2_nw[2][1]),
    .cast_ready_o_2_1                              (cast_ready_nw_2_pe[2][1]),
    .merge_data_i_2_1                              (merge_data_pe_2_nw[2][1]),
    .merge_valid_i_2_1                             (merge_valid_pe_2_nw[2][1]),
    .merge_ready_o_2_1                             (merge_ready_nw_2_pe[2][1]),
    .gather_data_i_2_1                             (gather_data_pe_2_nw[2][1]),
    .gather_valid_i_2_1                            (gather_valid_pe_2_nw[2][1]),
    .gather_ready_o_2_1                            (gather_ready_nw_2_pe[2][1]),

    .cast_data_o_2_1                               (cast_data_nw_2_pe[2][1]),
    .cast_valid_o_2_1                              (cast_valid_nw_2_pe[2][1]),
    .cast_ready_i_2_1                              (cast_ready_pe_2_nw[2][1]),
    .merge_data_o_2_1                              (merge_data_nw_2_pe[2][1]),
    .merge_valid_o_2_1                             (merge_valid_nw_2_pe[2][1]),
    .merge_ready_i_2_1                             (merge_ready_pe_2_nw[2][1]),
    .gather_data_o_2_1                             (gather_data_nw_2_pe[2][1]),
    .gather_valid_o_2_1                            (gather_valid_nw_2_pe[2][1]),
    .gather_ready_i_2_1                            (gather_ready_pe_2_nw[2][1]),
    .cast_data_i_2_2                               (cast_data_pe_2_nw[2][2]),
    .cast_valid_i_2_2                              (cast_valid_pe_2_nw[2][2]),
    .cast_ready_o_2_2                              (cast_ready_nw_2_pe[2][2]),
    .merge_data_i_2_2                              (merge_data_pe_2_nw[2][2]),
    .merge_valid_i_2_2                             (merge_valid_pe_2_nw[2][2]),
    .merge_ready_o_2_2                             (merge_ready_nw_2_pe[2][2]),
    .gather_data_i_2_2                             (gather_data_pe_2_nw[2][2]),
    .gather_valid_i_2_2                            (gather_valid_pe_2_nw[2][2]),
    .gather_ready_o_2_2                            (gather_ready_nw_2_pe[2][2]),

    .cast_data_o_2_2                               (cast_data_nw_2_pe[2][2]),
    .cast_valid_o_2_2                              (cast_valid_nw_2_pe[2][2]),
    .cast_ready_i_2_2                              (cast_ready_pe_2_nw[2][2]),
    .merge_data_o_2_2                              (merge_data_nw_2_pe[2][2]),
    .merge_valid_o_2_2                             (merge_valid_nw_2_pe[2][2]),
    .merge_ready_i_2_2                             (merge_ready_pe_2_nw[2][2]),
    .gather_data_o_2_2                             (gather_data_nw_2_pe[2][2]),
    .gather_valid_o_2_2                            (gather_valid_nw_2_pe[2][2]),
    .gather_ready_i_2_2                            (gather_ready_pe_2_nw[2][2]),
    .cast_data_i_2_3                               (cast_data_pe_2_nw[2][3]),
    .cast_valid_i_2_3                              (cast_valid_pe_2_nw[2][3]),
    .cast_ready_o_2_3                              (cast_ready_nw_2_pe[2][3]),
    .merge_data_i_2_3                              (merge_data_pe_2_nw[2][3]),
    .merge_valid_i_2_3                             (merge_valid_pe_2_nw[2][3]),
    .merge_ready_o_2_3                             (merge_ready_nw_2_pe[2][3]),
    .gather_data_i_2_3                             (gather_data_pe_2_nw[2][3]),
    .gather_valid_i_2_3                            (gather_valid_pe_2_nw[2][3]),
    .gather_ready_o_2_3                            (gather_ready_nw_2_pe[2][3]),

    .cast_data_o_2_3                               (cast_data_nw_2_pe[2][3]),
    .cast_valid_o_2_3                              (cast_valid_nw_2_pe[2][3]),
    .cast_ready_i_2_3                              (cast_ready_pe_2_nw[2][3]),
    .merge_data_o_2_3                              (merge_data_nw_2_pe[2][3]),
    .merge_valid_o_2_3                             (merge_valid_nw_2_pe[2][3]),
    .merge_ready_i_2_3                             (merge_ready_pe_2_nw[2][3]),
    .gather_data_o_2_3                             (gather_data_nw_2_pe[2][3]),
    .gather_valid_o_2_3                            (gather_valid_nw_2_pe[2][3]),
    .gather_ready_i_2_3                            (gather_ready_pe_2_nw[2][3]),
    .cast_data_i_2_4                               (cast_data_pe_2_nw[2][4]),
    .cast_valid_i_2_4                              (cast_valid_pe_2_nw[2][4]),
    .cast_ready_o_2_4                              (cast_ready_nw_2_pe[2][4]),
    .merge_data_i_2_4                              (merge_data_pe_2_nw[2][4]),
    .merge_valid_i_2_4                             (merge_valid_pe_2_nw[2][4]),
    .merge_ready_o_2_4                             (merge_ready_nw_2_pe[2][4]),
    .gather_data_i_2_4                             (gather_data_pe_2_nw[2][4]),
    .gather_valid_i_2_4                            (gather_valid_pe_2_nw[2][4]),
    .gather_ready_o_2_4                            (gather_ready_nw_2_pe[2][4]),

    .cast_data_o_2_4                               (cast_data_nw_2_pe[2][4]),
    .cast_valid_o_2_4                              (cast_valid_nw_2_pe[2][4]),
    .cast_ready_i_2_4                              (cast_ready_pe_2_nw[2][4]),
    .merge_data_o_2_4                              (merge_data_nw_2_pe[2][4]),
    .merge_valid_o_2_4                             (merge_valid_nw_2_pe[2][4]),
    .merge_ready_i_2_4                             (merge_ready_pe_2_nw[2][4]),
    .gather_data_o_2_4                             (gather_data_nw_2_pe[2][4]),
    .gather_valid_o_2_4                            (gather_valid_nw_2_pe[2][4]),
    .gather_ready_i_2_4                            (gather_ready_pe_2_nw[2][4]),
    .cast_data_i_2_5                               (cast_data_pe_2_nw[2][5]),
    .cast_valid_i_2_5                              (cast_valid_pe_2_nw[2][5]),
    .cast_ready_o_2_5                              (cast_ready_nw_2_pe[2][5]),
    .merge_data_i_2_5                              (merge_data_pe_2_nw[2][5]),
    .merge_valid_i_2_5                             (merge_valid_pe_2_nw[2][5]),
    .merge_ready_o_2_5                             (merge_ready_nw_2_pe[2][5]),
    .gather_data_i_2_5                             (gather_data_pe_2_nw[2][5]),
    .gather_valid_i_2_5                            (gather_valid_pe_2_nw[2][5]),
    .gather_ready_o_2_5                            (gather_ready_nw_2_pe[2][5]),

    .cast_data_o_2_5                               (cast_data_nw_2_pe[2][5]),
    .cast_valid_o_2_5                              (cast_valid_nw_2_pe[2][5]),
    .cast_ready_i_2_5                              (cast_ready_pe_2_nw[2][5]),
    .merge_data_o_2_5                              (merge_data_nw_2_pe[2][5]),
    .merge_valid_o_2_5                             (merge_valid_nw_2_pe[2][5]),
    .merge_ready_i_2_5                             (merge_ready_pe_2_nw[2][5]),
    .gather_data_o_2_5                             (gather_data_nw_2_pe[2][5]),
    .gather_valid_o_2_5                            (gather_valid_nw_2_pe[2][5]),
    .gather_ready_i_2_5                            (gather_ready_pe_2_nw[2][5]),
    .cast_data_i_2_6                               (cast_data_pe_2_nw[2][6]),
    .cast_valid_i_2_6                              (cast_valid_pe_2_nw[2][6]),
    .cast_ready_o_2_6                              (cast_ready_nw_2_pe[2][6]),
    .merge_data_i_2_6                              (merge_data_pe_2_nw[2][6]),
    .merge_valid_i_2_6                             (merge_valid_pe_2_nw[2][6]),
    .merge_ready_o_2_6                             (merge_ready_nw_2_pe[2][6]),
    .gather_data_i_2_6                             (gather_data_pe_2_nw[2][6]),
    .gather_valid_i_2_6                            (gather_valid_pe_2_nw[2][6]),
    .gather_ready_o_2_6                            (gather_ready_nw_2_pe[2][6]),

    .cast_data_o_2_6                               (cast_data_nw_2_pe[2][6]),
    .cast_valid_o_2_6                              (cast_valid_nw_2_pe[2][6]),
    .cast_ready_i_2_6                              (cast_ready_pe_2_nw[2][6]),
    .merge_data_o_2_6                              (merge_data_nw_2_pe[2][6]),
    .merge_valid_o_2_6                             (merge_valid_nw_2_pe[2][6]),
    .merge_ready_i_2_6                             (merge_ready_pe_2_nw[2][6]),
    .gather_data_o_2_6                             (gather_data_nw_2_pe[2][6]),
    .gather_valid_o_2_6                            (gather_valid_nw_2_pe[2][6]),
    .gather_ready_i_2_6                            (gather_ready_pe_2_nw[2][6]),
    .cast_data_i_2_7                               (cast_data_pe_2_nw[2][7]),
    .cast_valid_i_2_7                              (cast_valid_pe_2_nw[2][7]),
    .cast_ready_o_2_7                              (cast_ready_nw_2_pe[2][7]),
    .merge_data_i_2_7                              (merge_data_pe_2_nw[2][7]),
    .merge_valid_i_2_7                             (merge_valid_pe_2_nw[2][7]),
    .merge_ready_o_2_7                             (merge_ready_nw_2_pe[2][7]),
    .gather_data_i_2_7                             (gather_data_pe_2_nw[2][7]),
    .gather_valid_i_2_7                            (gather_valid_pe_2_nw[2][7]),
    .gather_ready_o_2_7                            (gather_ready_nw_2_pe[2][7]),

    .cast_data_o_2_7                               (cast_data_nw_2_pe[2][7]),
    .cast_valid_o_2_7                              (cast_valid_nw_2_pe[2][7]),
    .cast_ready_i_2_7                              (cast_ready_pe_2_nw[2][7]),
    .merge_data_o_2_7                              (merge_data_nw_2_pe[2][7]),
    .merge_valid_o_2_7                             (merge_valid_nw_2_pe[2][7]),
    .merge_ready_i_2_7                             (merge_ready_pe_2_nw[2][7]),
    .gather_data_o_2_7                             (gather_data_nw_2_pe[2][7]),
    .gather_valid_o_2_7                            (gather_valid_nw_2_pe[2][7]),
    .gather_ready_i_2_7                            (gather_ready_pe_2_nw[2][7]),
    .cast_data_i_2_8                               (cast_data_pe_2_nw[2][8]),
    .cast_valid_i_2_8                              (cast_valid_pe_2_nw[2][8]),
    .cast_ready_o_2_8                              (cast_ready_nw_2_pe[2][8]),
    .merge_data_i_2_8                              (merge_data_pe_2_nw[2][8]),
    .merge_valid_i_2_8                             (merge_valid_pe_2_nw[2][8]),
    .merge_ready_o_2_8                             (merge_ready_nw_2_pe[2][8]),
    .gather_data_i_2_8                             (gather_data_pe_2_nw[2][8]),
    .gather_valid_i_2_8                            (gather_valid_pe_2_nw[2][8]),
    .gather_ready_o_2_8                            (gather_ready_nw_2_pe[2][8]),

    .cast_data_o_2_8                               (cast_data_nw_2_pe[2][8]),
    .cast_valid_o_2_8                              (cast_valid_nw_2_pe[2][8]),
    .cast_ready_i_2_8                              (cast_ready_pe_2_nw[2][8]),
    .merge_data_o_2_8                              (merge_data_nw_2_pe[2][8]),
    .merge_valid_o_2_8                             (merge_valid_nw_2_pe[2][8]),
    .merge_ready_i_2_8                             (merge_ready_pe_2_nw[2][8]),
    .gather_data_o_2_8                             (gather_data_nw_2_pe[2][8]),
    .gather_valid_o_2_8                            (gather_valid_nw_2_pe[2][8]),
    .gather_ready_i_2_8                            (gather_ready_pe_2_nw[2][8]),
    .cast_data_i_2_9                               (cast_data_pe_2_nw[2][9]),
    .cast_valid_i_2_9                              (cast_valid_pe_2_nw[2][9]),
    .cast_ready_o_2_9                              (cast_ready_nw_2_pe[2][9]),
    .merge_data_i_2_9                              (merge_data_pe_2_nw[2][9]),
    .merge_valid_i_2_9                             (merge_valid_pe_2_nw[2][9]),
    .merge_ready_o_2_9                             (merge_ready_nw_2_pe[2][9]),
    .gather_data_i_2_9                             (gather_data_pe_2_nw[2][9]),
    .gather_valid_i_2_9                            (gather_valid_pe_2_nw[2][9]),
    .gather_ready_o_2_9                            (gather_ready_nw_2_pe[2][9]),

    .cast_data_o_2_9                               (cast_data_nw_2_pe[2][9]),
    .cast_valid_o_2_9                              (cast_valid_nw_2_pe[2][9]),
    .cast_ready_i_2_9                              (cast_ready_pe_2_nw[2][9]),
    .merge_data_o_2_9                              (merge_data_nw_2_pe[2][9]),
    .merge_valid_o_2_9                             (merge_valid_nw_2_pe[2][9]),
    .merge_ready_i_2_9                             (merge_ready_pe_2_nw[2][9]),
    .gather_data_o_2_9                             (gather_data_nw_2_pe[2][9]),
    .gather_valid_o_2_9                            (gather_valid_nw_2_pe[2][9]),
    .gather_ready_i_2_9                            (gather_ready_pe_2_nw[2][9]),
    .cast_data_i_2_10                               (cast_data_pe_2_nw[2][10]),
    .cast_valid_i_2_10                              (cast_valid_pe_2_nw[2][10]),
    .cast_ready_o_2_10                              (cast_ready_nw_2_pe[2][10]),
    .merge_data_i_2_10                              (merge_data_pe_2_nw[2][10]),
    .merge_valid_i_2_10                             (merge_valid_pe_2_nw[2][10]),
    .merge_ready_o_2_10                             (merge_ready_nw_2_pe[2][10]),
    .gather_data_i_2_10                             (gather_data_pe_2_nw[2][10]),
    .gather_valid_i_2_10                            (gather_valid_pe_2_nw[2][10]),
    .gather_ready_o_2_10                            (gather_ready_nw_2_pe[2][10]),

    .cast_data_o_2_10                               (cast_data_nw_2_pe[2][10]),
    .cast_valid_o_2_10                              (cast_valid_nw_2_pe[2][10]),
    .cast_ready_i_2_10                              (cast_ready_pe_2_nw[2][10]),
    .merge_data_o_2_10                              (merge_data_nw_2_pe[2][10]),
    .merge_valid_o_2_10                             (merge_valid_nw_2_pe[2][10]),
    .merge_ready_i_2_10                             (merge_ready_pe_2_nw[2][10]),
    .gather_data_o_2_10                             (gather_data_nw_2_pe[2][10]),
    .gather_valid_o_2_10                            (gather_valid_nw_2_pe[2][10]),
    .gather_ready_i_2_10                            (gather_ready_pe_2_nw[2][10]),
    .cast_data_i_2_11                               (cast_data_pe_2_nw[2][11]),
    .cast_valid_i_2_11                              (cast_valid_pe_2_nw[2][11]),
    .cast_ready_o_2_11                              (cast_ready_nw_2_pe[2][11]),
    .merge_data_i_2_11                              (merge_data_pe_2_nw[2][11]),
    .merge_valid_i_2_11                             (merge_valid_pe_2_nw[2][11]),
    .merge_ready_o_2_11                             (merge_ready_nw_2_pe[2][11]),
    .gather_data_i_2_11                             (gather_data_pe_2_nw[2][11]),
    .gather_valid_i_2_11                            (gather_valid_pe_2_nw[2][11]),
    .gather_ready_o_2_11                            (gather_ready_nw_2_pe[2][11]),

    .cast_data_o_2_11                               (cast_data_nw_2_pe[2][11]),
    .cast_valid_o_2_11                              (cast_valid_nw_2_pe[2][11]),
    .cast_ready_i_2_11                              (cast_ready_pe_2_nw[2][11]),
    .merge_data_o_2_11                              (merge_data_nw_2_pe[2][11]),
    .merge_valid_o_2_11                             (merge_valid_nw_2_pe[2][11]),
    .merge_ready_i_2_11                             (merge_ready_pe_2_nw[2][11]),
    .gather_data_o_2_11                             (gather_data_nw_2_pe[2][11]),
    .gather_valid_o_2_11                            (gather_valid_nw_2_pe[2][11]),
    .gather_ready_i_2_11                            (gather_ready_pe_2_nw[2][11]),
    .cast_data_i_2_12                               (cast_data_pe_2_nw[2][12]),
    .cast_valid_i_2_12                              (cast_valid_pe_2_nw[2][12]),
    .cast_ready_o_2_12                              (cast_ready_nw_2_pe[2][12]),
    .merge_data_i_2_12                              (merge_data_pe_2_nw[2][12]),
    .merge_valid_i_2_12                             (merge_valid_pe_2_nw[2][12]),
    .merge_ready_o_2_12                             (merge_ready_nw_2_pe[2][12]),
    .gather_data_i_2_12                             (gather_data_pe_2_nw[2][12]),
    .gather_valid_i_2_12                            (gather_valid_pe_2_nw[2][12]),
    .gather_ready_o_2_12                            (gather_ready_nw_2_pe[2][12]),

    .cast_data_o_2_12                               (cast_data_nw_2_pe[2][12]),
    .cast_valid_o_2_12                              (cast_valid_nw_2_pe[2][12]),
    .cast_ready_i_2_12                              (cast_ready_pe_2_nw[2][12]),
    .merge_data_o_2_12                              (merge_data_nw_2_pe[2][12]),
    .merge_valid_o_2_12                             (merge_valid_nw_2_pe[2][12]),
    .merge_ready_i_2_12                             (merge_ready_pe_2_nw[2][12]),
    .gather_data_o_2_12                             (gather_data_nw_2_pe[2][12]),
    .gather_valid_o_2_12                            (gather_valid_nw_2_pe[2][12]),
    .gather_ready_i_2_12                            (gather_ready_pe_2_nw[2][12]),
    .cast_data_i_2_13                               (cast_data_pe_2_nw[2][13]),
    .cast_valid_i_2_13                              (cast_valid_pe_2_nw[2][13]),
    .cast_ready_o_2_13                              (cast_ready_nw_2_pe[2][13]),
    .merge_data_i_2_13                              (merge_data_pe_2_nw[2][13]),
    .merge_valid_i_2_13                             (merge_valid_pe_2_nw[2][13]),
    .merge_ready_o_2_13                             (merge_ready_nw_2_pe[2][13]),
    .gather_data_i_2_13                             (gather_data_pe_2_nw[2][13]),
    .gather_valid_i_2_13                            (gather_valid_pe_2_nw[2][13]),
    .gather_ready_o_2_13                            (gather_ready_nw_2_pe[2][13]),

    .cast_data_o_2_13                               (cast_data_nw_2_pe[2][13]),
    .cast_valid_o_2_13                              (cast_valid_nw_2_pe[2][13]),
    .cast_ready_i_2_13                              (cast_ready_pe_2_nw[2][13]),
    .merge_data_o_2_13                              (merge_data_nw_2_pe[2][13]),
    .merge_valid_o_2_13                             (merge_valid_nw_2_pe[2][13]),
    .merge_ready_i_2_13                             (merge_ready_pe_2_nw[2][13]),
    .gather_data_o_2_13                             (gather_data_nw_2_pe[2][13]),
    .gather_valid_o_2_13                            (gather_valid_nw_2_pe[2][13]),
    .gather_ready_i_2_13                            (gather_ready_pe_2_nw[2][13]),
    .cast_data_i_2_14                               (cast_data_pe_2_nw[2][14]),
    .cast_valid_i_2_14                              (cast_valid_pe_2_nw[2][14]),
    .cast_ready_o_2_14                              (cast_ready_nw_2_pe[2][14]),
    .merge_data_i_2_14                              (merge_data_pe_2_nw[2][14]),
    .merge_valid_i_2_14                             (merge_valid_pe_2_nw[2][14]),
    .merge_ready_o_2_14                             (merge_ready_nw_2_pe[2][14]),
    .gather_data_i_2_14                             (gather_data_pe_2_nw[2][14]),
    .gather_valid_i_2_14                            (gather_valid_pe_2_nw[2][14]),
    .gather_ready_o_2_14                            (gather_ready_nw_2_pe[2][14]),

    .cast_data_o_2_14                               (cast_data_nw_2_pe[2][14]),
    .cast_valid_o_2_14                              (cast_valid_nw_2_pe[2][14]),
    .cast_ready_i_2_14                              (cast_ready_pe_2_nw[2][14]),
    .merge_data_o_2_14                              (merge_data_nw_2_pe[2][14]),
    .merge_valid_o_2_14                             (merge_valid_nw_2_pe[2][14]),
    .merge_ready_i_2_14                             (merge_ready_pe_2_nw[2][14]),
    .gather_data_o_2_14                             (gather_data_nw_2_pe[2][14]),
    .gather_valid_o_2_14                            (gather_valid_nw_2_pe[2][14]),
    .gather_ready_i_2_14                            (gather_ready_pe_2_nw[2][14]),
    .cast_data_i_2_15                               (cast_data_pe_2_nw[2][15]),
    .cast_valid_i_2_15                              (cast_valid_pe_2_nw[2][15]),
    .cast_ready_o_2_15                              (cast_ready_nw_2_pe[2][15]),
    .merge_data_i_2_15                              (merge_data_pe_2_nw[2][15]),
    .merge_valid_i_2_15                             (merge_valid_pe_2_nw[2][15]),
    .merge_ready_o_2_15                             (merge_ready_nw_2_pe[2][15]),
    .gather_data_i_2_15                             (gather_data_pe_2_nw[2][15]),
    .gather_valid_i_2_15                            (gather_valid_pe_2_nw[2][15]),
    .gather_ready_o_2_15                            (gather_ready_nw_2_pe[2][15]),

    .cast_data_o_2_15                               (cast_data_nw_2_pe[2][15]),
    .cast_valid_o_2_15                              (cast_valid_nw_2_pe[2][15]),
    .cast_ready_i_2_15                              (cast_ready_pe_2_nw[2][15]),
    .merge_data_o_2_15                              (merge_data_nw_2_pe[2][15]),
    .merge_valid_o_2_15                             (merge_valid_nw_2_pe[2][15]),
    .merge_ready_i_2_15                             (merge_ready_pe_2_nw[2][15]),
    .gather_data_o_2_15                             (gather_data_nw_2_pe[2][15]),
    .gather_valid_o_2_15                            (gather_valid_nw_2_pe[2][15]),
    .gather_ready_i_2_15                            (gather_ready_pe_2_nw[2][15]),
    .cast_data_i_2_16                               (cast_data_pe_2_nw[2][16]),
    .cast_valid_i_2_16                              (cast_valid_pe_2_nw[2][16]),
    .cast_ready_o_2_16                              (cast_ready_nw_2_pe[2][16]),
    .merge_data_i_2_16                              (merge_data_pe_2_nw[2][16]),
    .merge_valid_i_2_16                             (merge_valid_pe_2_nw[2][16]),
    .merge_ready_o_2_16                             (merge_ready_nw_2_pe[2][16]),
    .gather_data_i_2_16                             (gather_data_pe_2_nw[2][16]),
    .gather_valid_i_2_16                            (gather_valid_pe_2_nw[2][16]),
    .gather_ready_o_2_16                            (gather_ready_nw_2_pe[2][16]),

    .cast_data_o_2_16                               (cast_data_nw_2_pe[2][16]),
    .cast_valid_o_2_16                              (cast_valid_nw_2_pe[2][16]),
    .cast_ready_i_2_16                              (cast_ready_pe_2_nw[2][16]),
    .merge_data_o_2_16                              (merge_data_nw_2_pe[2][16]),
    .merge_valid_o_2_16                             (merge_valid_nw_2_pe[2][16]),
    .merge_ready_i_2_16                             (merge_ready_pe_2_nw[2][16]),
    .gather_data_o_2_16                             (gather_data_nw_2_pe[2][16]),
    .gather_valid_o_2_16                            (gather_valid_nw_2_pe[2][16]),
    .gather_ready_i_2_16                            (gather_ready_pe_2_nw[2][16]),
    .cast_data_i_2_17                               (cast_data_pe_2_nw[2][17]),
    .cast_valid_i_2_17                              (cast_valid_pe_2_nw[2][17]),
    .cast_ready_o_2_17                              (cast_ready_nw_2_pe[2][17]),
    .merge_data_i_2_17                              (merge_data_pe_2_nw[2][17]),
    .merge_valid_i_2_17                             (merge_valid_pe_2_nw[2][17]),
    .merge_ready_o_2_17                             (merge_ready_nw_2_pe[2][17]),
    .gather_data_i_2_17                             (gather_data_pe_2_nw[2][17]),
    .gather_valid_i_2_17                            (gather_valid_pe_2_nw[2][17]),
    .gather_ready_o_2_17                            (gather_ready_nw_2_pe[2][17]),

    .cast_data_o_2_17                               (cast_data_nw_2_pe[2][17]),
    .cast_valid_o_2_17                              (cast_valid_nw_2_pe[2][17]),
    .cast_ready_i_2_17                              (cast_ready_pe_2_nw[2][17]),
    .merge_data_o_2_17                              (merge_data_nw_2_pe[2][17]),
    .merge_valid_o_2_17                             (merge_valid_nw_2_pe[2][17]),
    .merge_ready_i_2_17                             (merge_ready_pe_2_nw[2][17]),
    .gather_data_o_2_17                             (gather_data_nw_2_pe[2][17]),
    .gather_valid_o_2_17                            (gather_valid_nw_2_pe[2][17]),
    .gather_ready_i_2_17                            (gather_ready_pe_2_nw[2][17]),
    .cast_data_i_2_18                               (cast_data_pe_2_nw[2][18]),
    .cast_valid_i_2_18                              (cast_valid_pe_2_nw[2][18]),
    .cast_ready_o_2_18                              (cast_ready_nw_2_pe[2][18]),
    .merge_data_i_2_18                              (merge_data_pe_2_nw[2][18]),
    .merge_valid_i_2_18                             (merge_valid_pe_2_nw[2][18]),
    .merge_ready_o_2_18                             (merge_ready_nw_2_pe[2][18]),
    .gather_data_i_2_18                             (gather_data_pe_2_nw[2][18]),
    .gather_valid_i_2_18                            (gather_valid_pe_2_nw[2][18]),
    .gather_ready_o_2_18                            (gather_ready_nw_2_pe[2][18]),

    .cast_data_o_2_18                               (cast_data_nw_2_pe[2][18]),
    .cast_valid_o_2_18                              (cast_valid_nw_2_pe[2][18]),
    .cast_ready_i_2_18                              (cast_ready_pe_2_nw[2][18]),
    .merge_data_o_2_18                              (merge_data_nw_2_pe[2][18]),
    .merge_valid_o_2_18                             (merge_valid_nw_2_pe[2][18]),
    .merge_ready_i_2_18                             (merge_ready_pe_2_nw[2][18]),
    .gather_data_o_2_18                             (gather_data_nw_2_pe[2][18]),
    .gather_valid_o_2_18                            (gather_valid_nw_2_pe[2][18]),
    .gather_ready_i_2_18                            (gather_ready_pe_2_nw[2][18]),
    .cast_data_i_2_19                               (cast_data_pe_2_nw[2][19]),
    .cast_valid_i_2_19                              (cast_valid_pe_2_nw[2][19]),
    .cast_ready_o_2_19                              (cast_ready_nw_2_pe[2][19]),
    .merge_data_i_2_19                              (merge_data_pe_2_nw[2][19]),
    .merge_valid_i_2_19                             (merge_valid_pe_2_nw[2][19]),
    .merge_ready_o_2_19                             (merge_ready_nw_2_pe[2][19]),
    .gather_data_i_2_19                             (gather_data_pe_2_nw[2][19]),
    .gather_valid_i_2_19                            (gather_valid_pe_2_nw[2][19]),
    .gather_ready_o_2_19                            (gather_ready_nw_2_pe[2][19]),

    .cast_data_o_2_19                               (cast_data_nw_2_pe[2][19]),
    .cast_valid_o_2_19                              (cast_valid_nw_2_pe[2][19]),
    .cast_ready_i_2_19                              (cast_ready_pe_2_nw[2][19]),
    .merge_data_o_2_19                              (merge_data_nw_2_pe[2][19]),
    .merge_valid_o_2_19                             (merge_valid_nw_2_pe[2][19]),
    .merge_ready_i_2_19                             (merge_ready_pe_2_nw[2][19]),
    .gather_data_o_2_19                             (gather_data_nw_2_pe[2][19]),
    .gather_valid_o_2_19                            (gather_valid_nw_2_pe[2][19]),
    .gather_ready_i_2_19                            (gather_ready_pe_2_nw[2][19]),
    .cast_data_i_2_20                               (cast_data_pe_2_nw[2][20]),
    .cast_valid_i_2_20                              (cast_valid_pe_2_nw[2][20]),
    .cast_ready_o_2_20                              (cast_ready_nw_2_pe[2][20]),
    .merge_data_i_2_20                              (merge_data_pe_2_nw[2][20]),
    .merge_valid_i_2_20                             (merge_valid_pe_2_nw[2][20]),
    .merge_ready_o_2_20                             (merge_ready_nw_2_pe[2][20]),
    .gather_data_i_2_20                             (gather_data_pe_2_nw[2][20]),
    .gather_valid_i_2_20                            (gather_valid_pe_2_nw[2][20]),
    .gather_ready_o_2_20                            (gather_ready_nw_2_pe[2][20]),

    .cast_data_o_2_20                               (cast_data_nw_2_pe[2][20]),
    .cast_valid_o_2_20                              (cast_valid_nw_2_pe[2][20]),
    .cast_ready_i_2_20                              (cast_ready_pe_2_nw[2][20]),
    .merge_data_o_2_20                              (merge_data_nw_2_pe[2][20]),
    .merge_valid_o_2_20                             (merge_valid_nw_2_pe[2][20]),
    .merge_ready_i_2_20                             (merge_ready_pe_2_nw[2][20]),
    .gather_data_o_2_20                             (gather_data_nw_2_pe[2][20]),
    .gather_valid_o_2_20                            (gather_valid_nw_2_pe[2][20]),
    .gather_ready_i_2_20                            (gather_ready_pe_2_nw[2][20]),
    .cast_data_i_2_21                               (cast_data_pe_2_nw[2][21]),
    .cast_valid_i_2_21                              (cast_valid_pe_2_nw[2][21]),
    .cast_ready_o_2_21                              (cast_ready_nw_2_pe[2][21]),
    .merge_data_i_2_21                              (merge_data_pe_2_nw[2][21]),
    .merge_valid_i_2_21                             (merge_valid_pe_2_nw[2][21]),
    .merge_ready_o_2_21                             (merge_ready_nw_2_pe[2][21]),
    .gather_data_i_2_21                             (gather_data_pe_2_nw[2][21]),
    .gather_valid_i_2_21                            (gather_valid_pe_2_nw[2][21]),
    .gather_ready_o_2_21                            (gather_ready_nw_2_pe[2][21]),

    .cast_data_o_2_21                               (cast_data_nw_2_pe[2][21]),
    .cast_valid_o_2_21                              (cast_valid_nw_2_pe[2][21]),
    .cast_ready_i_2_21                              (cast_ready_pe_2_nw[2][21]),
    .merge_data_o_2_21                              (merge_data_nw_2_pe[2][21]),
    .merge_valid_o_2_21                             (merge_valid_nw_2_pe[2][21]),
    .merge_ready_i_2_21                             (merge_ready_pe_2_nw[2][21]),
    .gather_data_o_2_21                             (gather_data_nw_2_pe[2][21]),
    .gather_valid_o_2_21                            (gather_valid_nw_2_pe[2][21]),
    .gather_ready_i_2_21                            (gather_ready_pe_2_nw[2][21]),
    .cast_data_i_2_22                               (cast_data_pe_2_nw[2][22]),
    .cast_valid_i_2_22                              (cast_valid_pe_2_nw[2][22]),
    .cast_ready_o_2_22                              (cast_ready_nw_2_pe[2][22]),
    .merge_data_i_2_22                              (merge_data_pe_2_nw[2][22]),
    .merge_valid_i_2_22                             (merge_valid_pe_2_nw[2][22]),
    .merge_ready_o_2_22                             (merge_ready_nw_2_pe[2][22]),
    .gather_data_i_2_22                             (gather_data_pe_2_nw[2][22]),
    .gather_valid_i_2_22                            (gather_valid_pe_2_nw[2][22]),
    .gather_ready_o_2_22                            (gather_ready_nw_2_pe[2][22]),

    .cast_data_o_2_22                               (cast_data_nw_2_pe[2][22]),
    .cast_valid_o_2_22                              (cast_valid_nw_2_pe[2][22]),
    .cast_ready_i_2_22                              (cast_ready_pe_2_nw[2][22]),
    .merge_data_o_2_22                              (merge_data_nw_2_pe[2][22]),
    .merge_valid_o_2_22                             (merge_valid_nw_2_pe[2][22]),
    .merge_ready_i_2_22                             (merge_ready_pe_2_nw[2][22]),
    .gather_data_o_2_22                             (gather_data_nw_2_pe[2][22]),
    .gather_valid_o_2_22                            (gather_valid_nw_2_pe[2][22]),
    .gather_ready_i_2_22                            (gather_ready_pe_2_nw[2][22]),
    .cast_data_i_2_23                               (cast_data_pe_2_nw[2][23]),
    .cast_valid_i_2_23                              (cast_valid_pe_2_nw[2][23]),
    .cast_ready_o_2_23                              (cast_ready_nw_2_pe[2][23]),
    .merge_data_i_2_23                              (merge_data_pe_2_nw[2][23]),
    .merge_valid_i_2_23                             (merge_valid_pe_2_nw[2][23]),
    .merge_ready_o_2_23                             (merge_ready_nw_2_pe[2][23]),
    .gather_data_i_2_23                             (gather_data_pe_2_nw[2][23]),
    .gather_valid_i_2_23                            (gather_valid_pe_2_nw[2][23]),
    .gather_ready_o_2_23                            (gather_ready_nw_2_pe[2][23]),

    .cast_data_o_2_23                               (cast_data_nw_2_pe[2][23]),
    .cast_valid_o_2_23                              (cast_valid_nw_2_pe[2][23]),
    .cast_ready_i_2_23                              (cast_ready_pe_2_nw[2][23]),
    .merge_data_o_2_23                              (merge_data_nw_2_pe[2][23]),
    .merge_valid_o_2_23                             (merge_valid_nw_2_pe[2][23]),
    .merge_ready_i_2_23                             (merge_ready_pe_2_nw[2][23]),
    .gather_data_o_2_23                             (gather_data_nw_2_pe[2][23]),
    .gather_valid_o_2_23                            (gather_valid_nw_2_pe[2][23]),
    .gather_ready_i_2_23                            (gather_ready_pe_2_nw[2][23]),
    .cast_data_i_2_24                               (cast_data_pe_2_nw[2][24]),
    .cast_valid_i_2_24                              (cast_valid_pe_2_nw[2][24]),
    .cast_ready_o_2_24                              (cast_ready_nw_2_pe[2][24]),
    .merge_data_i_2_24                              (merge_data_pe_2_nw[2][24]),
    .merge_valid_i_2_24                             (merge_valid_pe_2_nw[2][24]),
    .merge_ready_o_2_24                             (merge_ready_nw_2_pe[2][24]),
    .gather_data_i_2_24                             (gather_data_pe_2_nw[2][24]),
    .gather_valid_i_2_24                            (gather_valid_pe_2_nw[2][24]),
    .gather_ready_o_2_24                            (gather_ready_nw_2_pe[2][24]),

    .cast_data_o_2_24                               (cast_data_nw_2_pe[2][24]),
    .cast_valid_o_2_24                              (cast_valid_nw_2_pe[2][24]),
    .cast_ready_i_2_24                              (cast_ready_pe_2_nw[2][24]),
    .merge_data_o_2_24                              (merge_data_nw_2_pe[2][24]),
    .merge_valid_o_2_24                             (merge_valid_nw_2_pe[2][24]),
    .merge_ready_i_2_24                             (merge_ready_pe_2_nw[2][24]),
    .gather_data_o_2_24                             (gather_data_nw_2_pe[2][24]),
    .gather_valid_o_2_24                            (gather_valid_nw_2_pe[2][24]),
    .gather_ready_i_2_24                            (gather_ready_pe_2_nw[2][24]),
    .cast_data_i_3_0                               (cast_data_pe_2_nw[3][0]),
    .cast_valid_i_3_0                              (cast_valid_pe_2_nw[3][0]),
    .cast_ready_o_3_0                              (cast_ready_nw_2_pe[3][0]),
    .merge_data_i_3_0                              (merge_data_pe_2_nw[3][0]),
    .merge_valid_i_3_0                             (merge_valid_pe_2_nw[3][0]),
    .merge_ready_o_3_0                             (merge_ready_nw_2_pe[3][0]),
    .gather_data_i_3_0                             (gather_data_pe_2_nw[3][0]),
    .gather_valid_i_3_0                            (gather_valid_pe_2_nw[3][0]),
    .gather_ready_o_3_0                            (gather_ready_nw_2_pe[3][0]),

    .cast_data_o_3_0                               (cast_data_nw_2_pe[3][0]),
    .cast_valid_o_3_0                              (cast_valid_nw_2_pe[3][0]),
    .cast_ready_i_3_0                              (cast_ready_pe_2_nw[3][0]),
    .merge_data_o_3_0                              (merge_data_nw_2_pe[3][0]),
    .merge_valid_o_3_0                             (merge_valid_nw_2_pe[3][0]),
    .merge_ready_i_3_0                             (merge_ready_pe_2_nw[3][0]),
    .gather_data_o_3_0                             (gather_data_nw_2_pe[3][0]),
    .gather_valid_o_3_0                            (gather_valid_nw_2_pe[3][0]),
    .gather_ready_i_3_0                            (gather_ready_pe_2_nw[3][0]),
    .cast_data_i_3_1                               (cast_data_pe_2_nw[3][1]),
    .cast_valid_i_3_1                              (cast_valid_pe_2_nw[3][1]),
    .cast_ready_o_3_1                              (cast_ready_nw_2_pe[3][1]),
    .merge_data_i_3_1                              (merge_data_pe_2_nw[3][1]),
    .merge_valid_i_3_1                             (merge_valid_pe_2_nw[3][1]),
    .merge_ready_o_3_1                             (merge_ready_nw_2_pe[3][1]),
    .gather_data_i_3_1                             (gather_data_pe_2_nw[3][1]),
    .gather_valid_i_3_1                            (gather_valid_pe_2_nw[3][1]),
    .gather_ready_o_3_1                            (gather_ready_nw_2_pe[3][1]),

    .cast_data_o_3_1                               (cast_data_nw_2_pe[3][1]),
    .cast_valid_o_3_1                              (cast_valid_nw_2_pe[3][1]),
    .cast_ready_i_3_1                              (cast_ready_pe_2_nw[3][1]),
    .merge_data_o_3_1                              (merge_data_nw_2_pe[3][1]),
    .merge_valid_o_3_1                             (merge_valid_nw_2_pe[3][1]),
    .merge_ready_i_3_1                             (merge_ready_pe_2_nw[3][1]),
    .gather_data_o_3_1                             (gather_data_nw_2_pe[3][1]),
    .gather_valid_o_3_1                            (gather_valid_nw_2_pe[3][1]),
    .gather_ready_i_3_1                            (gather_ready_pe_2_nw[3][1]),
    .cast_data_i_3_2                               (cast_data_pe_2_nw[3][2]),
    .cast_valid_i_3_2                              (cast_valid_pe_2_nw[3][2]),
    .cast_ready_o_3_2                              (cast_ready_nw_2_pe[3][2]),
    .merge_data_i_3_2                              (merge_data_pe_2_nw[3][2]),
    .merge_valid_i_3_2                             (merge_valid_pe_2_nw[3][2]),
    .merge_ready_o_3_2                             (merge_ready_nw_2_pe[3][2]),
    .gather_data_i_3_2                             (gather_data_pe_2_nw[3][2]),
    .gather_valid_i_3_2                            (gather_valid_pe_2_nw[3][2]),
    .gather_ready_o_3_2                            (gather_ready_nw_2_pe[3][2]),

    .cast_data_o_3_2                               (cast_data_nw_2_pe[3][2]),
    .cast_valid_o_3_2                              (cast_valid_nw_2_pe[3][2]),
    .cast_ready_i_3_2                              (cast_ready_pe_2_nw[3][2]),
    .merge_data_o_3_2                              (merge_data_nw_2_pe[3][2]),
    .merge_valid_o_3_2                             (merge_valid_nw_2_pe[3][2]),
    .merge_ready_i_3_2                             (merge_ready_pe_2_nw[3][2]),
    .gather_data_o_3_2                             (gather_data_nw_2_pe[3][2]),
    .gather_valid_o_3_2                            (gather_valid_nw_2_pe[3][2]),
    .gather_ready_i_3_2                            (gather_ready_pe_2_nw[3][2]),
    .cast_data_i_3_3                               (cast_data_pe_2_nw[3][3]),
    .cast_valid_i_3_3                              (cast_valid_pe_2_nw[3][3]),
    .cast_ready_o_3_3                              (cast_ready_nw_2_pe[3][3]),
    .merge_data_i_3_3                              (merge_data_pe_2_nw[3][3]),
    .merge_valid_i_3_3                             (merge_valid_pe_2_nw[3][3]),
    .merge_ready_o_3_3                             (merge_ready_nw_2_pe[3][3]),
    .gather_data_i_3_3                             (gather_data_pe_2_nw[3][3]),
    .gather_valid_i_3_3                            (gather_valid_pe_2_nw[3][3]),
    .gather_ready_o_3_3                            (gather_ready_nw_2_pe[3][3]),

    .cast_data_o_3_3                               (cast_data_nw_2_pe[3][3]),
    .cast_valid_o_3_3                              (cast_valid_nw_2_pe[3][3]),
    .cast_ready_i_3_3                              (cast_ready_pe_2_nw[3][3]),
    .merge_data_o_3_3                              (merge_data_nw_2_pe[3][3]),
    .merge_valid_o_3_3                             (merge_valid_nw_2_pe[3][3]),
    .merge_ready_i_3_3                             (merge_ready_pe_2_nw[3][3]),
    .gather_data_o_3_3                             (gather_data_nw_2_pe[3][3]),
    .gather_valid_o_3_3                            (gather_valid_nw_2_pe[3][3]),
    .gather_ready_i_3_3                            (gather_ready_pe_2_nw[3][3]),
    .cast_data_i_3_4                               (cast_data_pe_2_nw[3][4]),
    .cast_valid_i_3_4                              (cast_valid_pe_2_nw[3][4]),
    .cast_ready_o_3_4                              (cast_ready_nw_2_pe[3][4]),
    .merge_data_i_3_4                              (merge_data_pe_2_nw[3][4]),
    .merge_valid_i_3_4                             (merge_valid_pe_2_nw[3][4]),
    .merge_ready_o_3_4                             (merge_ready_nw_2_pe[3][4]),
    .gather_data_i_3_4                             (gather_data_pe_2_nw[3][4]),
    .gather_valid_i_3_4                            (gather_valid_pe_2_nw[3][4]),
    .gather_ready_o_3_4                            (gather_ready_nw_2_pe[3][4]),

    .cast_data_o_3_4                               (cast_data_nw_2_pe[3][4]),
    .cast_valid_o_3_4                              (cast_valid_nw_2_pe[3][4]),
    .cast_ready_i_3_4                              (cast_ready_pe_2_nw[3][4]),
    .merge_data_o_3_4                              (merge_data_nw_2_pe[3][4]),
    .merge_valid_o_3_4                             (merge_valid_nw_2_pe[3][4]),
    .merge_ready_i_3_4                             (merge_ready_pe_2_nw[3][4]),
    .gather_data_o_3_4                             (gather_data_nw_2_pe[3][4]),
    .gather_valid_o_3_4                            (gather_valid_nw_2_pe[3][4]),
    .gather_ready_i_3_4                            (gather_ready_pe_2_nw[3][4]),
    .cast_data_i_3_5                               (cast_data_pe_2_nw[3][5]),
    .cast_valid_i_3_5                              (cast_valid_pe_2_nw[3][5]),
    .cast_ready_o_3_5                              (cast_ready_nw_2_pe[3][5]),
    .merge_data_i_3_5                              (merge_data_pe_2_nw[3][5]),
    .merge_valid_i_3_5                             (merge_valid_pe_2_nw[3][5]),
    .merge_ready_o_3_5                             (merge_ready_nw_2_pe[3][5]),
    .gather_data_i_3_5                             (gather_data_pe_2_nw[3][5]),
    .gather_valid_i_3_5                            (gather_valid_pe_2_nw[3][5]),
    .gather_ready_o_3_5                            (gather_ready_nw_2_pe[3][5]),

    .cast_data_o_3_5                               (cast_data_nw_2_pe[3][5]),
    .cast_valid_o_3_5                              (cast_valid_nw_2_pe[3][5]),
    .cast_ready_i_3_5                              (cast_ready_pe_2_nw[3][5]),
    .merge_data_o_3_5                              (merge_data_nw_2_pe[3][5]),
    .merge_valid_o_3_5                             (merge_valid_nw_2_pe[3][5]),
    .merge_ready_i_3_5                             (merge_ready_pe_2_nw[3][5]),
    .gather_data_o_3_5                             (gather_data_nw_2_pe[3][5]),
    .gather_valid_o_3_5                            (gather_valid_nw_2_pe[3][5]),
    .gather_ready_i_3_5                            (gather_ready_pe_2_nw[3][5]),
    .cast_data_i_3_6                               (cast_data_pe_2_nw[3][6]),
    .cast_valid_i_3_6                              (cast_valid_pe_2_nw[3][6]),
    .cast_ready_o_3_6                              (cast_ready_nw_2_pe[3][6]),
    .merge_data_i_3_6                              (merge_data_pe_2_nw[3][6]),
    .merge_valid_i_3_6                             (merge_valid_pe_2_nw[3][6]),
    .merge_ready_o_3_6                             (merge_ready_nw_2_pe[3][6]),
    .gather_data_i_3_6                             (gather_data_pe_2_nw[3][6]),
    .gather_valid_i_3_6                            (gather_valid_pe_2_nw[3][6]),
    .gather_ready_o_3_6                            (gather_ready_nw_2_pe[3][6]),

    .cast_data_o_3_6                               (cast_data_nw_2_pe[3][6]),
    .cast_valid_o_3_6                              (cast_valid_nw_2_pe[3][6]),
    .cast_ready_i_3_6                              (cast_ready_pe_2_nw[3][6]),
    .merge_data_o_3_6                              (merge_data_nw_2_pe[3][6]),
    .merge_valid_o_3_6                             (merge_valid_nw_2_pe[3][6]),
    .merge_ready_i_3_6                             (merge_ready_pe_2_nw[3][6]),
    .gather_data_o_3_6                             (gather_data_nw_2_pe[3][6]),
    .gather_valid_o_3_6                            (gather_valid_nw_2_pe[3][6]),
    .gather_ready_i_3_6                            (gather_ready_pe_2_nw[3][6]),
    .cast_data_i_3_7                               (cast_data_pe_2_nw[3][7]),
    .cast_valid_i_3_7                              (cast_valid_pe_2_nw[3][7]),
    .cast_ready_o_3_7                              (cast_ready_nw_2_pe[3][7]),
    .merge_data_i_3_7                              (merge_data_pe_2_nw[3][7]),
    .merge_valid_i_3_7                             (merge_valid_pe_2_nw[3][7]),
    .merge_ready_o_3_7                             (merge_ready_nw_2_pe[3][7]),
    .gather_data_i_3_7                             (gather_data_pe_2_nw[3][7]),
    .gather_valid_i_3_7                            (gather_valid_pe_2_nw[3][7]),
    .gather_ready_o_3_7                            (gather_ready_nw_2_pe[3][7]),

    .cast_data_o_3_7                               (cast_data_nw_2_pe[3][7]),
    .cast_valid_o_3_7                              (cast_valid_nw_2_pe[3][7]),
    .cast_ready_i_3_7                              (cast_ready_pe_2_nw[3][7]),
    .merge_data_o_3_7                              (merge_data_nw_2_pe[3][7]),
    .merge_valid_o_3_7                             (merge_valid_nw_2_pe[3][7]),
    .merge_ready_i_3_7                             (merge_ready_pe_2_nw[3][7]),
    .gather_data_o_3_7                             (gather_data_nw_2_pe[3][7]),
    .gather_valid_o_3_7                            (gather_valid_nw_2_pe[3][7]),
    .gather_ready_i_3_7                            (gather_ready_pe_2_nw[3][7]),
    .cast_data_i_3_8                               (cast_data_pe_2_nw[3][8]),
    .cast_valid_i_3_8                              (cast_valid_pe_2_nw[3][8]),
    .cast_ready_o_3_8                              (cast_ready_nw_2_pe[3][8]),
    .merge_data_i_3_8                              (merge_data_pe_2_nw[3][8]),
    .merge_valid_i_3_8                             (merge_valid_pe_2_nw[3][8]),
    .merge_ready_o_3_8                             (merge_ready_nw_2_pe[3][8]),
    .gather_data_i_3_8                             (gather_data_pe_2_nw[3][8]),
    .gather_valid_i_3_8                            (gather_valid_pe_2_nw[3][8]),
    .gather_ready_o_3_8                            (gather_ready_nw_2_pe[3][8]),

    .cast_data_o_3_8                               (cast_data_nw_2_pe[3][8]),
    .cast_valid_o_3_8                              (cast_valid_nw_2_pe[3][8]),
    .cast_ready_i_3_8                              (cast_ready_pe_2_nw[3][8]),
    .merge_data_o_3_8                              (merge_data_nw_2_pe[3][8]),
    .merge_valid_o_3_8                             (merge_valid_nw_2_pe[3][8]),
    .merge_ready_i_3_8                             (merge_ready_pe_2_nw[3][8]),
    .gather_data_o_3_8                             (gather_data_nw_2_pe[3][8]),
    .gather_valid_o_3_8                            (gather_valid_nw_2_pe[3][8]),
    .gather_ready_i_3_8                            (gather_ready_pe_2_nw[3][8]),
    .cast_data_i_3_9                               (cast_data_pe_2_nw[3][9]),
    .cast_valid_i_3_9                              (cast_valid_pe_2_nw[3][9]),
    .cast_ready_o_3_9                              (cast_ready_nw_2_pe[3][9]),
    .merge_data_i_3_9                              (merge_data_pe_2_nw[3][9]),
    .merge_valid_i_3_9                             (merge_valid_pe_2_nw[3][9]),
    .merge_ready_o_3_9                             (merge_ready_nw_2_pe[3][9]),
    .gather_data_i_3_9                             (gather_data_pe_2_nw[3][9]),
    .gather_valid_i_3_9                            (gather_valid_pe_2_nw[3][9]),
    .gather_ready_o_3_9                            (gather_ready_nw_2_pe[3][9]),

    .cast_data_o_3_9                               (cast_data_nw_2_pe[3][9]),
    .cast_valid_o_3_9                              (cast_valid_nw_2_pe[3][9]),
    .cast_ready_i_3_9                              (cast_ready_pe_2_nw[3][9]),
    .merge_data_o_3_9                              (merge_data_nw_2_pe[3][9]),
    .merge_valid_o_3_9                             (merge_valid_nw_2_pe[3][9]),
    .merge_ready_i_3_9                             (merge_ready_pe_2_nw[3][9]),
    .gather_data_o_3_9                             (gather_data_nw_2_pe[3][9]),
    .gather_valid_o_3_9                            (gather_valid_nw_2_pe[3][9]),
    .gather_ready_i_3_9                            (gather_ready_pe_2_nw[3][9]),
    .cast_data_i_3_10                               (cast_data_pe_2_nw[3][10]),
    .cast_valid_i_3_10                              (cast_valid_pe_2_nw[3][10]),
    .cast_ready_o_3_10                              (cast_ready_nw_2_pe[3][10]),
    .merge_data_i_3_10                              (merge_data_pe_2_nw[3][10]),
    .merge_valid_i_3_10                             (merge_valid_pe_2_nw[3][10]),
    .merge_ready_o_3_10                             (merge_ready_nw_2_pe[3][10]),
    .gather_data_i_3_10                             (gather_data_pe_2_nw[3][10]),
    .gather_valid_i_3_10                            (gather_valid_pe_2_nw[3][10]),
    .gather_ready_o_3_10                            (gather_ready_nw_2_pe[3][10]),

    .cast_data_o_3_10                               (cast_data_nw_2_pe[3][10]),
    .cast_valid_o_3_10                              (cast_valid_nw_2_pe[3][10]),
    .cast_ready_i_3_10                              (cast_ready_pe_2_nw[3][10]),
    .merge_data_o_3_10                              (merge_data_nw_2_pe[3][10]),
    .merge_valid_o_3_10                             (merge_valid_nw_2_pe[3][10]),
    .merge_ready_i_3_10                             (merge_ready_pe_2_nw[3][10]),
    .gather_data_o_3_10                             (gather_data_nw_2_pe[3][10]),
    .gather_valid_o_3_10                            (gather_valid_nw_2_pe[3][10]),
    .gather_ready_i_3_10                            (gather_ready_pe_2_nw[3][10]),
    .cast_data_i_3_11                               (cast_data_pe_2_nw[3][11]),
    .cast_valid_i_3_11                              (cast_valid_pe_2_nw[3][11]),
    .cast_ready_o_3_11                              (cast_ready_nw_2_pe[3][11]),
    .merge_data_i_3_11                              (merge_data_pe_2_nw[3][11]),
    .merge_valid_i_3_11                             (merge_valid_pe_2_nw[3][11]),
    .merge_ready_o_3_11                             (merge_ready_nw_2_pe[3][11]),
    .gather_data_i_3_11                             (gather_data_pe_2_nw[3][11]),
    .gather_valid_i_3_11                            (gather_valid_pe_2_nw[3][11]),
    .gather_ready_o_3_11                            (gather_ready_nw_2_pe[3][11]),

    .cast_data_o_3_11                               (cast_data_nw_2_pe[3][11]),
    .cast_valid_o_3_11                              (cast_valid_nw_2_pe[3][11]),
    .cast_ready_i_3_11                              (cast_ready_pe_2_nw[3][11]),
    .merge_data_o_3_11                              (merge_data_nw_2_pe[3][11]),
    .merge_valid_o_3_11                             (merge_valid_nw_2_pe[3][11]),
    .merge_ready_i_3_11                             (merge_ready_pe_2_nw[3][11]),
    .gather_data_o_3_11                             (gather_data_nw_2_pe[3][11]),
    .gather_valid_o_3_11                            (gather_valid_nw_2_pe[3][11]),
    .gather_ready_i_3_11                            (gather_ready_pe_2_nw[3][11]),
    .cast_data_i_3_12                               (cast_data_pe_2_nw[3][12]),
    .cast_valid_i_3_12                              (cast_valid_pe_2_nw[3][12]),
    .cast_ready_o_3_12                              (cast_ready_nw_2_pe[3][12]),
    .merge_data_i_3_12                              (merge_data_pe_2_nw[3][12]),
    .merge_valid_i_3_12                             (merge_valid_pe_2_nw[3][12]),
    .merge_ready_o_3_12                             (merge_ready_nw_2_pe[3][12]),
    .gather_data_i_3_12                             (gather_data_pe_2_nw[3][12]),
    .gather_valid_i_3_12                            (gather_valid_pe_2_nw[3][12]),
    .gather_ready_o_3_12                            (gather_ready_nw_2_pe[3][12]),

    .cast_data_o_3_12                               (cast_data_nw_2_pe[3][12]),
    .cast_valid_o_3_12                              (cast_valid_nw_2_pe[3][12]),
    .cast_ready_i_3_12                              (cast_ready_pe_2_nw[3][12]),
    .merge_data_o_3_12                              (merge_data_nw_2_pe[3][12]),
    .merge_valid_o_3_12                             (merge_valid_nw_2_pe[3][12]),
    .merge_ready_i_3_12                             (merge_ready_pe_2_nw[3][12]),
    .gather_data_o_3_12                             (gather_data_nw_2_pe[3][12]),
    .gather_valid_o_3_12                            (gather_valid_nw_2_pe[3][12]),
    .gather_ready_i_3_12                            (gather_ready_pe_2_nw[3][12]),
    .cast_data_i_3_13                               (cast_data_pe_2_nw[3][13]),
    .cast_valid_i_3_13                              (cast_valid_pe_2_nw[3][13]),
    .cast_ready_o_3_13                              (cast_ready_nw_2_pe[3][13]),
    .merge_data_i_3_13                              (merge_data_pe_2_nw[3][13]),
    .merge_valid_i_3_13                             (merge_valid_pe_2_nw[3][13]),
    .merge_ready_o_3_13                             (merge_ready_nw_2_pe[3][13]),
    .gather_data_i_3_13                             (gather_data_pe_2_nw[3][13]),
    .gather_valid_i_3_13                            (gather_valid_pe_2_nw[3][13]),
    .gather_ready_o_3_13                            (gather_ready_nw_2_pe[3][13]),

    .cast_data_o_3_13                               (cast_data_nw_2_pe[3][13]),
    .cast_valid_o_3_13                              (cast_valid_nw_2_pe[3][13]),
    .cast_ready_i_3_13                              (cast_ready_pe_2_nw[3][13]),
    .merge_data_o_3_13                              (merge_data_nw_2_pe[3][13]),
    .merge_valid_o_3_13                             (merge_valid_nw_2_pe[3][13]),
    .merge_ready_i_3_13                             (merge_ready_pe_2_nw[3][13]),
    .gather_data_o_3_13                             (gather_data_nw_2_pe[3][13]),
    .gather_valid_o_3_13                            (gather_valid_nw_2_pe[3][13]),
    .gather_ready_i_3_13                            (gather_ready_pe_2_nw[3][13]),
    .cast_data_i_3_14                               (cast_data_pe_2_nw[3][14]),
    .cast_valid_i_3_14                              (cast_valid_pe_2_nw[3][14]),
    .cast_ready_o_3_14                              (cast_ready_nw_2_pe[3][14]),
    .merge_data_i_3_14                              (merge_data_pe_2_nw[3][14]),
    .merge_valid_i_3_14                             (merge_valid_pe_2_nw[3][14]),
    .merge_ready_o_3_14                             (merge_ready_nw_2_pe[3][14]),
    .gather_data_i_3_14                             (gather_data_pe_2_nw[3][14]),
    .gather_valid_i_3_14                            (gather_valid_pe_2_nw[3][14]),
    .gather_ready_o_3_14                            (gather_ready_nw_2_pe[3][14]),

    .cast_data_o_3_14                               (cast_data_nw_2_pe[3][14]),
    .cast_valid_o_3_14                              (cast_valid_nw_2_pe[3][14]),
    .cast_ready_i_3_14                              (cast_ready_pe_2_nw[3][14]),
    .merge_data_o_3_14                              (merge_data_nw_2_pe[3][14]),
    .merge_valid_o_3_14                             (merge_valid_nw_2_pe[3][14]),
    .merge_ready_i_3_14                             (merge_ready_pe_2_nw[3][14]),
    .gather_data_o_3_14                             (gather_data_nw_2_pe[3][14]),
    .gather_valid_o_3_14                            (gather_valid_nw_2_pe[3][14]),
    .gather_ready_i_3_14                            (gather_ready_pe_2_nw[3][14]),
    .cast_data_i_3_15                               (cast_data_pe_2_nw[3][15]),
    .cast_valid_i_3_15                              (cast_valid_pe_2_nw[3][15]),
    .cast_ready_o_3_15                              (cast_ready_nw_2_pe[3][15]),
    .merge_data_i_3_15                              (merge_data_pe_2_nw[3][15]),
    .merge_valid_i_3_15                             (merge_valid_pe_2_nw[3][15]),
    .merge_ready_o_3_15                             (merge_ready_nw_2_pe[3][15]),
    .gather_data_i_3_15                             (gather_data_pe_2_nw[3][15]),
    .gather_valid_i_3_15                            (gather_valid_pe_2_nw[3][15]),
    .gather_ready_o_3_15                            (gather_ready_nw_2_pe[3][15]),

    .cast_data_o_3_15                               (cast_data_nw_2_pe[3][15]),
    .cast_valid_o_3_15                              (cast_valid_nw_2_pe[3][15]),
    .cast_ready_i_3_15                              (cast_ready_pe_2_nw[3][15]),
    .merge_data_o_3_15                              (merge_data_nw_2_pe[3][15]),
    .merge_valid_o_3_15                             (merge_valid_nw_2_pe[3][15]),
    .merge_ready_i_3_15                             (merge_ready_pe_2_nw[3][15]),
    .gather_data_o_3_15                             (gather_data_nw_2_pe[3][15]),
    .gather_valid_o_3_15                            (gather_valid_nw_2_pe[3][15]),
    .gather_ready_i_3_15                            (gather_ready_pe_2_nw[3][15]),
    .cast_data_i_3_16                               (cast_data_pe_2_nw[3][16]),
    .cast_valid_i_3_16                              (cast_valid_pe_2_nw[3][16]),
    .cast_ready_o_3_16                              (cast_ready_nw_2_pe[3][16]),
    .merge_data_i_3_16                              (merge_data_pe_2_nw[3][16]),
    .merge_valid_i_3_16                             (merge_valid_pe_2_nw[3][16]),
    .merge_ready_o_3_16                             (merge_ready_nw_2_pe[3][16]),
    .gather_data_i_3_16                             (gather_data_pe_2_nw[3][16]),
    .gather_valid_i_3_16                            (gather_valid_pe_2_nw[3][16]),
    .gather_ready_o_3_16                            (gather_ready_nw_2_pe[3][16]),

    .cast_data_o_3_16                               (cast_data_nw_2_pe[3][16]),
    .cast_valid_o_3_16                              (cast_valid_nw_2_pe[3][16]),
    .cast_ready_i_3_16                              (cast_ready_pe_2_nw[3][16]),
    .merge_data_o_3_16                              (merge_data_nw_2_pe[3][16]),
    .merge_valid_o_3_16                             (merge_valid_nw_2_pe[3][16]),
    .merge_ready_i_3_16                             (merge_ready_pe_2_nw[3][16]),
    .gather_data_o_3_16                             (gather_data_nw_2_pe[3][16]),
    .gather_valid_o_3_16                            (gather_valid_nw_2_pe[3][16]),
    .gather_ready_i_3_16                            (gather_ready_pe_2_nw[3][16]),
    .cast_data_i_3_17                               (cast_data_pe_2_nw[3][17]),
    .cast_valid_i_3_17                              (cast_valid_pe_2_nw[3][17]),
    .cast_ready_o_3_17                              (cast_ready_nw_2_pe[3][17]),
    .merge_data_i_3_17                              (merge_data_pe_2_nw[3][17]),
    .merge_valid_i_3_17                             (merge_valid_pe_2_nw[3][17]),
    .merge_ready_o_3_17                             (merge_ready_nw_2_pe[3][17]),
    .gather_data_i_3_17                             (gather_data_pe_2_nw[3][17]),
    .gather_valid_i_3_17                            (gather_valid_pe_2_nw[3][17]),
    .gather_ready_o_3_17                            (gather_ready_nw_2_pe[3][17]),

    .cast_data_o_3_17                               (cast_data_nw_2_pe[3][17]),
    .cast_valid_o_3_17                              (cast_valid_nw_2_pe[3][17]),
    .cast_ready_i_3_17                              (cast_ready_pe_2_nw[3][17]),
    .merge_data_o_3_17                              (merge_data_nw_2_pe[3][17]),
    .merge_valid_o_3_17                             (merge_valid_nw_2_pe[3][17]),
    .merge_ready_i_3_17                             (merge_ready_pe_2_nw[3][17]),
    .gather_data_o_3_17                             (gather_data_nw_2_pe[3][17]),
    .gather_valid_o_3_17                            (gather_valid_nw_2_pe[3][17]),
    .gather_ready_i_3_17                            (gather_ready_pe_2_nw[3][17]),
    .cast_data_i_3_18                               (cast_data_pe_2_nw[3][18]),
    .cast_valid_i_3_18                              (cast_valid_pe_2_nw[3][18]),
    .cast_ready_o_3_18                              (cast_ready_nw_2_pe[3][18]),
    .merge_data_i_3_18                              (merge_data_pe_2_nw[3][18]),
    .merge_valid_i_3_18                             (merge_valid_pe_2_nw[3][18]),
    .merge_ready_o_3_18                             (merge_ready_nw_2_pe[3][18]),
    .gather_data_i_3_18                             (gather_data_pe_2_nw[3][18]),
    .gather_valid_i_3_18                            (gather_valid_pe_2_nw[3][18]),
    .gather_ready_o_3_18                            (gather_ready_nw_2_pe[3][18]),

    .cast_data_o_3_18                               (cast_data_nw_2_pe[3][18]),
    .cast_valid_o_3_18                              (cast_valid_nw_2_pe[3][18]),
    .cast_ready_i_3_18                              (cast_ready_pe_2_nw[3][18]),
    .merge_data_o_3_18                              (merge_data_nw_2_pe[3][18]),
    .merge_valid_o_3_18                             (merge_valid_nw_2_pe[3][18]),
    .merge_ready_i_3_18                             (merge_ready_pe_2_nw[3][18]),
    .gather_data_o_3_18                             (gather_data_nw_2_pe[3][18]),
    .gather_valid_o_3_18                            (gather_valid_nw_2_pe[3][18]),
    .gather_ready_i_3_18                            (gather_ready_pe_2_nw[3][18]),
    .cast_data_i_3_19                               (cast_data_pe_2_nw[3][19]),
    .cast_valid_i_3_19                              (cast_valid_pe_2_nw[3][19]),
    .cast_ready_o_3_19                              (cast_ready_nw_2_pe[3][19]),
    .merge_data_i_3_19                              (merge_data_pe_2_nw[3][19]),
    .merge_valid_i_3_19                             (merge_valid_pe_2_nw[3][19]),
    .merge_ready_o_3_19                             (merge_ready_nw_2_pe[3][19]),
    .gather_data_i_3_19                             (gather_data_pe_2_nw[3][19]),
    .gather_valid_i_3_19                            (gather_valid_pe_2_nw[3][19]),
    .gather_ready_o_3_19                            (gather_ready_nw_2_pe[3][19]),

    .cast_data_o_3_19                               (cast_data_nw_2_pe[3][19]),
    .cast_valid_o_3_19                              (cast_valid_nw_2_pe[3][19]),
    .cast_ready_i_3_19                              (cast_ready_pe_2_nw[3][19]),
    .merge_data_o_3_19                              (merge_data_nw_2_pe[3][19]),
    .merge_valid_o_3_19                             (merge_valid_nw_2_pe[3][19]),
    .merge_ready_i_3_19                             (merge_ready_pe_2_nw[3][19]),
    .gather_data_o_3_19                             (gather_data_nw_2_pe[3][19]),
    .gather_valid_o_3_19                            (gather_valid_nw_2_pe[3][19]),
    .gather_ready_i_3_19                            (gather_ready_pe_2_nw[3][19]),
    .cast_data_i_3_20                               (cast_data_pe_2_nw[3][20]),
    .cast_valid_i_3_20                              (cast_valid_pe_2_nw[3][20]),
    .cast_ready_o_3_20                              (cast_ready_nw_2_pe[3][20]),
    .merge_data_i_3_20                              (merge_data_pe_2_nw[3][20]),
    .merge_valid_i_3_20                             (merge_valid_pe_2_nw[3][20]),
    .merge_ready_o_3_20                             (merge_ready_nw_2_pe[3][20]),
    .gather_data_i_3_20                             (gather_data_pe_2_nw[3][20]),
    .gather_valid_i_3_20                            (gather_valid_pe_2_nw[3][20]),
    .gather_ready_o_3_20                            (gather_ready_nw_2_pe[3][20]),

    .cast_data_o_3_20                               (cast_data_nw_2_pe[3][20]),
    .cast_valid_o_3_20                              (cast_valid_nw_2_pe[3][20]),
    .cast_ready_i_3_20                              (cast_ready_pe_2_nw[3][20]),
    .merge_data_o_3_20                              (merge_data_nw_2_pe[3][20]),
    .merge_valid_o_3_20                             (merge_valid_nw_2_pe[3][20]),
    .merge_ready_i_3_20                             (merge_ready_pe_2_nw[3][20]),
    .gather_data_o_3_20                             (gather_data_nw_2_pe[3][20]),
    .gather_valid_o_3_20                            (gather_valid_nw_2_pe[3][20]),
    .gather_ready_i_3_20                            (gather_ready_pe_2_nw[3][20]),
    .cast_data_i_3_21                               (cast_data_pe_2_nw[3][21]),
    .cast_valid_i_3_21                              (cast_valid_pe_2_nw[3][21]),
    .cast_ready_o_3_21                              (cast_ready_nw_2_pe[3][21]),
    .merge_data_i_3_21                              (merge_data_pe_2_nw[3][21]),
    .merge_valid_i_3_21                             (merge_valid_pe_2_nw[3][21]),
    .merge_ready_o_3_21                             (merge_ready_nw_2_pe[3][21]),
    .gather_data_i_3_21                             (gather_data_pe_2_nw[3][21]),
    .gather_valid_i_3_21                            (gather_valid_pe_2_nw[3][21]),
    .gather_ready_o_3_21                            (gather_ready_nw_2_pe[3][21]),

    .cast_data_o_3_21                               (cast_data_nw_2_pe[3][21]),
    .cast_valid_o_3_21                              (cast_valid_nw_2_pe[3][21]),
    .cast_ready_i_3_21                              (cast_ready_pe_2_nw[3][21]),
    .merge_data_o_3_21                              (merge_data_nw_2_pe[3][21]),
    .merge_valid_o_3_21                             (merge_valid_nw_2_pe[3][21]),
    .merge_ready_i_3_21                             (merge_ready_pe_2_nw[3][21]),
    .gather_data_o_3_21                             (gather_data_nw_2_pe[3][21]),
    .gather_valid_o_3_21                            (gather_valid_nw_2_pe[3][21]),
    .gather_ready_i_3_21                            (gather_ready_pe_2_nw[3][21]),
    .cast_data_i_3_22                               (cast_data_pe_2_nw[3][22]),
    .cast_valid_i_3_22                              (cast_valid_pe_2_nw[3][22]),
    .cast_ready_o_3_22                              (cast_ready_nw_2_pe[3][22]),
    .merge_data_i_3_22                              (merge_data_pe_2_nw[3][22]),
    .merge_valid_i_3_22                             (merge_valid_pe_2_nw[3][22]),
    .merge_ready_o_3_22                             (merge_ready_nw_2_pe[3][22]),
    .gather_data_i_3_22                             (gather_data_pe_2_nw[3][22]),
    .gather_valid_i_3_22                            (gather_valid_pe_2_nw[3][22]),
    .gather_ready_o_3_22                            (gather_ready_nw_2_pe[3][22]),

    .cast_data_o_3_22                               (cast_data_nw_2_pe[3][22]),
    .cast_valid_o_3_22                              (cast_valid_nw_2_pe[3][22]),
    .cast_ready_i_3_22                              (cast_ready_pe_2_nw[3][22]),
    .merge_data_o_3_22                              (merge_data_nw_2_pe[3][22]),
    .merge_valid_o_3_22                             (merge_valid_nw_2_pe[3][22]),
    .merge_ready_i_3_22                             (merge_ready_pe_2_nw[3][22]),
    .gather_data_o_3_22                             (gather_data_nw_2_pe[3][22]),
    .gather_valid_o_3_22                            (gather_valid_nw_2_pe[3][22]),
    .gather_ready_i_3_22                            (gather_ready_pe_2_nw[3][22]),
    .cast_data_i_3_23                               (cast_data_pe_2_nw[3][23]),
    .cast_valid_i_3_23                              (cast_valid_pe_2_nw[3][23]),
    .cast_ready_o_3_23                              (cast_ready_nw_2_pe[3][23]),
    .merge_data_i_3_23                              (merge_data_pe_2_nw[3][23]),
    .merge_valid_i_3_23                             (merge_valid_pe_2_nw[3][23]),
    .merge_ready_o_3_23                             (merge_ready_nw_2_pe[3][23]),
    .gather_data_i_3_23                             (gather_data_pe_2_nw[3][23]),
    .gather_valid_i_3_23                            (gather_valid_pe_2_nw[3][23]),
    .gather_ready_o_3_23                            (gather_ready_nw_2_pe[3][23]),

    .cast_data_o_3_23                               (cast_data_nw_2_pe[3][23]),
    .cast_valid_o_3_23                              (cast_valid_nw_2_pe[3][23]),
    .cast_ready_i_3_23                              (cast_ready_pe_2_nw[3][23]),
    .merge_data_o_3_23                              (merge_data_nw_2_pe[3][23]),
    .merge_valid_o_3_23                             (merge_valid_nw_2_pe[3][23]),
    .merge_ready_i_3_23                             (merge_ready_pe_2_nw[3][23]),
    .gather_data_o_3_23                             (gather_data_nw_2_pe[3][23]),
    .gather_valid_o_3_23                            (gather_valid_nw_2_pe[3][23]),
    .gather_ready_i_3_23                            (gather_ready_pe_2_nw[3][23]),
    .cast_data_i_3_24                               (cast_data_pe_2_nw[3][24]),
    .cast_valid_i_3_24                              (cast_valid_pe_2_nw[3][24]),
    .cast_ready_o_3_24                              (cast_ready_nw_2_pe[3][24]),
    .merge_data_i_3_24                              (merge_data_pe_2_nw[3][24]),
    .merge_valid_i_3_24                             (merge_valid_pe_2_nw[3][24]),
    .merge_ready_o_3_24                             (merge_ready_nw_2_pe[3][24]),
    .gather_data_i_3_24                             (gather_data_pe_2_nw[3][24]),
    .gather_valid_i_3_24                            (gather_valid_pe_2_nw[3][24]),
    .gather_ready_o_3_24                            (gather_ready_nw_2_pe[3][24]),

    .cast_data_o_3_24                               (cast_data_nw_2_pe[3][24]),
    .cast_valid_o_3_24                              (cast_valid_nw_2_pe[3][24]),
    .cast_ready_i_3_24                              (cast_ready_pe_2_nw[3][24]),
    .merge_data_o_3_24                              (merge_data_nw_2_pe[3][24]),
    .merge_valid_o_3_24                             (merge_valid_nw_2_pe[3][24]),
    .merge_ready_i_3_24                             (merge_ready_pe_2_nw[3][24]),
    .gather_data_o_3_24                             (gather_data_nw_2_pe[3][24]),
    .gather_valid_o_3_24                            (gather_valid_nw_2_pe[3][24]),
    .gather_ready_i_3_24                            (gather_ready_pe_2_nw[3][24]),
    .cast_data_i_4_0                               (cast_data_pe_2_nw[4][0]),
    .cast_valid_i_4_0                              (cast_valid_pe_2_nw[4][0]),
    .cast_ready_o_4_0                              (cast_ready_nw_2_pe[4][0]),
    .merge_data_i_4_0                              (merge_data_pe_2_nw[4][0]),
    .merge_valid_i_4_0                             (merge_valid_pe_2_nw[4][0]),
    .merge_ready_o_4_0                             (merge_ready_nw_2_pe[4][0]),
    .gather_data_i_4_0                             (gather_data_pe_2_nw[4][0]),
    .gather_valid_i_4_0                            (gather_valid_pe_2_nw[4][0]),
    .gather_ready_o_4_0                            (gather_ready_nw_2_pe[4][0]),

    .cast_data_o_4_0                               (cast_data_nw_2_pe[4][0]),
    .cast_valid_o_4_0                              (cast_valid_nw_2_pe[4][0]),
    .cast_ready_i_4_0                              (cast_ready_pe_2_nw[4][0]),
    .merge_data_o_4_0                              (merge_data_nw_2_pe[4][0]),
    .merge_valid_o_4_0                             (merge_valid_nw_2_pe[4][0]),
    .merge_ready_i_4_0                             (merge_ready_pe_2_nw[4][0]),
    .gather_data_o_4_0                             (gather_data_nw_2_pe[4][0]),
    .gather_valid_o_4_0                            (gather_valid_nw_2_pe[4][0]),
    .gather_ready_i_4_0                            (gather_ready_pe_2_nw[4][0]),
    .cast_data_i_4_1                               (cast_data_pe_2_nw[4][1]),
    .cast_valid_i_4_1                              (cast_valid_pe_2_nw[4][1]),
    .cast_ready_o_4_1                              (cast_ready_nw_2_pe[4][1]),
    .merge_data_i_4_1                              (merge_data_pe_2_nw[4][1]),
    .merge_valid_i_4_1                             (merge_valid_pe_2_nw[4][1]),
    .merge_ready_o_4_1                             (merge_ready_nw_2_pe[4][1]),
    .gather_data_i_4_1                             (gather_data_pe_2_nw[4][1]),
    .gather_valid_i_4_1                            (gather_valid_pe_2_nw[4][1]),
    .gather_ready_o_4_1                            (gather_ready_nw_2_pe[4][1]),

    .cast_data_o_4_1                               (cast_data_nw_2_pe[4][1]),
    .cast_valid_o_4_1                              (cast_valid_nw_2_pe[4][1]),
    .cast_ready_i_4_1                              (cast_ready_pe_2_nw[4][1]),
    .merge_data_o_4_1                              (merge_data_nw_2_pe[4][1]),
    .merge_valid_o_4_1                             (merge_valid_nw_2_pe[4][1]),
    .merge_ready_i_4_1                             (merge_ready_pe_2_nw[4][1]),
    .gather_data_o_4_1                             (gather_data_nw_2_pe[4][1]),
    .gather_valid_o_4_1                            (gather_valid_nw_2_pe[4][1]),
    .gather_ready_i_4_1                            (gather_ready_pe_2_nw[4][1]),
    .cast_data_i_4_2                               (cast_data_pe_2_nw[4][2]),
    .cast_valid_i_4_2                              (cast_valid_pe_2_nw[4][2]),
    .cast_ready_o_4_2                              (cast_ready_nw_2_pe[4][2]),
    .merge_data_i_4_2                              (merge_data_pe_2_nw[4][2]),
    .merge_valid_i_4_2                             (merge_valid_pe_2_nw[4][2]),
    .merge_ready_o_4_2                             (merge_ready_nw_2_pe[4][2]),
    .gather_data_i_4_2                             (gather_data_pe_2_nw[4][2]),
    .gather_valid_i_4_2                            (gather_valid_pe_2_nw[4][2]),
    .gather_ready_o_4_2                            (gather_ready_nw_2_pe[4][2]),

    .cast_data_o_4_2                               (cast_data_nw_2_pe[4][2]),
    .cast_valid_o_4_2                              (cast_valid_nw_2_pe[4][2]),
    .cast_ready_i_4_2                              (cast_ready_pe_2_nw[4][2]),
    .merge_data_o_4_2                              (merge_data_nw_2_pe[4][2]),
    .merge_valid_o_4_2                             (merge_valid_nw_2_pe[4][2]),
    .merge_ready_i_4_2                             (merge_ready_pe_2_nw[4][2]),
    .gather_data_o_4_2                             (gather_data_nw_2_pe[4][2]),
    .gather_valid_o_4_2                            (gather_valid_nw_2_pe[4][2]),
    .gather_ready_i_4_2                            (gather_ready_pe_2_nw[4][2]),
    .cast_data_i_4_3                               (cast_data_pe_2_nw[4][3]),
    .cast_valid_i_4_3                              (cast_valid_pe_2_nw[4][3]),
    .cast_ready_o_4_3                              (cast_ready_nw_2_pe[4][3]),
    .merge_data_i_4_3                              (merge_data_pe_2_nw[4][3]),
    .merge_valid_i_4_3                             (merge_valid_pe_2_nw[4][3]),
    .merge_ready_o_4_3                             (merge_ready_nw_2_pe[4][3]),
    .gather_data_i_4_3                             (gather_data_pe_2_nw[4][3]),
    .gather_valid_i_4_3                            (gather_valid_pe_2_nw[4][3]),
    .gather_ready_o_4_3                            (gather_ready_nw_2_pe[4][3]),

    .cast_data_o_4_3                               (cast_data_nw_2_pe[4][3]),
    .cast_valid_o_4_3                              (cast_valid_nw_2_pe[4][3]),
    .cast_ready_i_4_3                              (cast_ready_pe_2_nw[4][3]),
    .merge_data_o_4_3                              (merge_data_nw_2_pe[4][3]),
    .merge_valid_o_4_3                             (merge_valid_nw_2_pe[4][3]),
    .merge_ready_i_4_3                             (merge_ready_pe_2_nw[4][3]),
    .gather_data_o_4_3                             (gather_data_nw_2_pe[4][3]),
    .gather_valid_o_4_3                            (gather_valid_nw_2_pe[4][3]),
    .gather_ready_i_4_3                            (gather_ready_pe_2_nw[4][3]),
    .cast_data_i_4_4                               (cast_data_pe_2_nw[4][4]),
    .cast_valid_i_4_4                              (cast_valid_pe_2_nw[4][4]),
    .cast_ready_o_4_4                              (cast_ready_nw_2_pe[4][4]),
    .merge_data_i_4_4                              (merge_data_pe_2_nw[4][4]),
    .merge_valid_i_4_4                             (merge_valid_pe_2_nw[4][4]),
    .merge_ready_o_4_4                             (merge_ready_nw_2_pe[4][4]),
    .gather_data_i_4_4                             (gather_data_pe_2_nw[4][4]),
    .gather_valid_i_4_4                            (gather_valid_pe_2_nw[4][4]),
    .gather_ready_o_4_4                            (gather_ready_nw_2_pe[4][4]),

    .cast_data_o_4_4                               (cast_data_nw_2_pe[4][4]),
    .cast_valid_o_4_4                              (cast_valid_nw_2_pe[4][4]),
    .cast_ready_i_4_4                              (cast_ready_pe_2_nw[4][4]),
    .merge_data_o_4_4                              (merge_data_nw_2_pe[4][4]),
    .merge_valid_o_4_4                             (merge_valid_nw_2_pe[4][4]),
    .merge_ready_i_4_4                             (merge_ready_pe_2_nw[4][4]),
    .gather_data_o_4_4                             (gather_data_nw_2_pe[4][4]),
    .gather_valid_o_4_4                            (gather_valid_nw_2_pe[4][4]),
    .gather_ready_i_4_4                            (gather_ready_pe_2_nw[4][4]),
    .cast_data_i_4_5                               (cast_data_pe_2_nw[4][5]),
    .cast_valid_i_4_5                              (cast_valid_pe_2_nw[4][5]),
    .cast_ready_o_4_5                              (cast_ready_nw_2_pe[4][5]),
    .merge_data_i_4_5                              (merge_data_pe_2_nw[4][5]),
    .merge_valid_i_4_5                             (merge_valid_pe_2_nw[4][5]),
    .merge_ready_o_4_5                             (merge_ready_nw_2_pe[4][5]),
    .gather_data_i_4_5                             (gather_data_pe_2_nw[4][5]),
    .gather_valid_i_4_5                            (gather_valid_pe_2_nw[4][5]),
    .gather_ready_o_4_5                            (gather_ready_nw_2_pe[4][5]),

    .cast_data_o_4_5                               (cast_data_nw_2_pe[4][5]),
    .cast_valid_o_4_5                              (cast_valid_nw_2_pe[4][5]),
    .cast_ready_i_4_5                              (cast_ready_pe_2_nw[4][5]),
    .merge_data_o_4_5                              (merge_data_nw_2_pe[4][5]),
    .merge_valid_o_4_5                             (merge_valid_nw_2_pe[4][5]),
    .merge_ready_i_4_5                             (merge_ready_pe_2_nw[4][5]),
    .gather_data_o_4_5                             (gather_data_nw_2_pe[4][5]),
    .gather_valid_o_4_5                            (gather_valid_nw_2_pe[4][5]),
    .gather_ready_i_4_5                            (gather_ready_pe_2_nw[4][5]),
    .cast_data_i_4_6                               (cast_data_pe_2_nw[4][6]),
    .cast_valid_i_4_6                              (cast_valid_pe_2_nw[4][6]),
    .cast_ready_o_4_6                              (cast_ready_nw_2_pe[4][6]),
    .merge_data_i_4_6                              (merge_data_pe_2_nw[4][6]),
    .merge_valid_i_4_6                             (merge_valid_pe_2_nw[4][6]),
    .merge_ready_o_4_6                             (merge_ready_nw_2_pe[4][6]),
    .gather_data_i_4_6                             (gather_data_pe_2_nw[4][6]),
    .gather_valid_i_4_6                            (gather_valid_pe_2_nw[4][6]),
    .gather_ready_o_4_6                            (gather_ready_nw_2_pe[4][6]),

    .cast_data_o_4_6                               (cast_data_nw_2_pe[4][6]),
    .cast_valid_o_4_6                              (cast_valid_nw_2_pe[4][6]),
    .cast_ready_i_4_6                              (cast_ready_pe_2_nw[4][6]),
    .merge_data_o_4_6                              (merge_data_nw_2_pe[4][6]),
    .merge_valid_o_4_6                             (merge_valid_nw_2_pe[4][6]),
    .merge_ready_i_4_6                             (merge_ready_pe_2_nw[4][6]),
    .gather_data_o_4_6                             (gather_data_nw_2_pe[4][6]),
    .gather_valid_o_4_6                            (gather_valid_nw_2_pe[4][6]),
    .gather_ready_i_4_6                            (gather_ready_pe_2_nw[4][6]),
    .cast_data_i_4_7                               (cast_data_pe_2_nw[4][7]),
    .cast_valid_i_4_7                              (cast_valid_pe_2_nw[4][7]),
    .cast_ready_o_4_7                              (cast_ready_nw_2_pe[4][7]),
    .merge_data_i_4_7                              (merge_data_pe_2_nw[4][7]),
    .merge_valid_i_4_7                             (merge_valid_pe_2_nw[4][7]),
    .merge_ready_o_4_7                             (merge_ready_nw_2_pe[4][7]),
    .gather_data_i_4_7                             (gather_data_pe_2_nw[4][7]),
    .gather_valid_i_4_7                            (gather_valid_pe_2_nw[4][7]),
    .gather_ready_o_4_7                            (gather_ready_nw_2_pe[4][7]),

    .cast_data_o_4_7                               (cast_data_nw_2_pe[4][7]),
    .cast_valid_o_4_7                              (cast_valid_nw_2_pe[4][7]),
    .cast_ready_i_4_7                              (cast_ready_pe_2_nw[4][7]),
    .merge_data_o_4_7                              (merge_data_nw_2_pe[4][7]),
    .merge_valid_o_4_7                             (merge_valid_nw_2_pe[4][7]),
    .merge_ready_i_4_7                             (merge_ready_pe_2_nw[4][7]),
    .gather_data_o_4_7                             (gather_data_nw_2_pe[4][7]),
    .gather_valid_o_4_7                            (gather_valid_nw_2_pe[4][7]),
    .gather_ready_i_4_7                            (gather_ready_pe_2_nw[4][7]),
    .cast_data_i_4_8                               (cast_data_pe_2_nw[4][8]),
    .cast_valid_i_4_8                              (cast_valid_pe_2_nw[4][8]),
    .cast_ready_o_4_8                              (cast_ready_nw_2_pe[4][8]),
    .merge_data_i_4_8                              (merge_data_pe_2_nw[4][8]),
    .merge_valid_i_4_8                             (merge_valid_pe_2_nw[4][8]),
    .merge_ready_o_4_8                             (merge_ready_nw_2_pe[4][8]),
    .gather_data_i_4_8                             (gather_data_pe_2_nw[4][8]),
    .gather_valid_i_4_8                            (gather_valid_pe_2_nw[4][8]),
    .gather_ready_o_4_8                            (gather_ready_nw_2_pe[4][8]),

    .cast_data_o_4_8                               (cast_data_nw_2_pe[4][8]),
    .cast_valid_o_4_8                              (cast_valid_nw_2_pe[4][8]),
    .cast_ready_i_4_8                              (cast_ready_pe_2_nw[4][8]),
    .merge_data_o_4_8                              (merge_data_nw_2_pe[4][8]),
    .merge_valid_o_4_8                             (merge_valid_nw_2_pe[4][8]),
    .merge_ready_i_4_8                             (merge_ready_pe_2_nw[4][8]),
    .gather_data_o_4_8                             (gather_data_nw_2_pe[4][8]),
    .gather_valid_o_4_8                            (gather_valid_nw_2_pe[4][8]),
    .gather_ready_i_4_8                            (gather_ready_pe_2_nw[4][8]),
    .cast_data_i_4_9                               (cast_data_pe_2_nw[4][9]),
    .cast_valid_i_4_9                              (cast_valid_pe_2_nw[4][9]),
    .cast_ready_o_4_9                              (cast_ready_nw_2_pe[4][9]),
    .merge_data_i_4_9                              (merge_data_pe_2_nw[4][9]),
    .merge_valid_i_4_9                             (merge_valid_pe_2_nw[4][9]),
    .merge_ready_o_4_9                             (merge_ready_nw_2_pe[4][9]),
    .gather_data_i_4_9                             (gather_data_pe_2_nw[4][9]),
    .gather_valid_i_4_9                            (gather_valid_pe_2_nw[4][9]),
    .gather_ready_o_4_9                            (gather_ready_nw_2_pe[4][9]),

    .cast_data_o_4_9                               (cast_data_nw_2_pe[4][9]),
    .cast_valid_o_4_9                              (cast_valid_nw_2_pe[4][9]),
    .cast_ready_i_4_9                              (cast_ready_pe_2_nw[4][9]),
    .merge_data_o_4_9                              (merge_data_nw_2_pe[4][9]),
    .merge_valid_o_4_9                             (merge_valid_nw_2_pe[4][9]),
    .merge_ready_i_4_9                             (merge_ready_pe_2_nw[4][9]),
    .gather_data_o_4_9                             (gather_data_nw_2_pe[4][9]),
    .gather_valid_o_4_9                            (gather_valid_nw_2_pe[4][9]),
    .gather_ready_i_4_9                            (gather_ready_pe_2_nw[4][9]),
    .cast_data_i_4_10                               (cast_data_pe_2_nw[4][10]),
    .cast_valid_i_4_10                              (cast_valid_pe_2_nw[4][10]),
    .cast_ready_o_4_10                              (cast_ready_nw_2_pe[4][10]),
    .merge_data_i_4_10                              (merge_data_pe_2_nw[4][10]),
    .merge_valid_i_4_10                             (merge_valid_pe_2_nw[4][10]),
    .merge_ready_o_4_10                             (merge_ready_nw_2_pe[4][10]),
    .gather_data_i_4_10                             (gather_data_pe_2_nw[4][10]),
    .gather_valid_i_4_10                            (gather_valid_pe_2_nw[4][10]),
    .gather_ready_o_4_10                            (gather_ready_nw_2_pe[4][10]),

    .cast_data_o_4_10                               (cast_data_nw_2_pe[4][10]),
    .cast_valid_o_4_10                              (cast_valid_nw_2_pe[4][10]),
    .cast_ready_i_4_10                              (cast_ready_pe_2_nw[4][10]),
    .merge_data_o_4_10                              (merge_data_nw_2_pe[4][10]),
    .merge_valid_o_4_10                             (merge_valid_nw_2_pe[4][10]),
    .merge_ready_i_4_10                             (merge_ready_pe_2_nw[4][10]),
    .gather_data_o_4_10                             (gather_data_nw_2_pe[4][10]),
    .gather_valid_o_4_10                            (gather_valid_nw_2_pe[4][10]),
    .gather_ready_i_4_10                            (gather_ready_pe_2_nw[4][10]),
    .cast_data_i_4_11                               (cast_data_pe_2_nw[4][11]),
    .cast_valid_i_4_11                              (cast_valid_pe_2_nw[4][11]),
    .cast_ready_o_4_11                              (cast_ready_nw_2_pe[4][11]),
    .merge_data_i_4_11                              (merge_data_pe_2_nw[4][11]),
    .merge_valid_i_4_11                             (merge_valid_pe_2_nw[4][11]),
    .merge_ready_o_4_11                             (merge_ready_nw_2_pe[4][11]),
    .gather_data_i_4_11                             (gather_data_pe_2_nw[4][11]),
    .gather_valid_i_4_11                            (gather_valid_pe_2_nw[4][11]),
    .gather_ready_o_4_11                            (gather_ready_nw_2_pe[4][11]),

    .cast_data_o_4_11                               (cast_data_nw_2_pe[4][11]),
    .cast_valid_o_4_11                              (cast_valid_nw_2_pe[4][11]),
    .cast_ready_i_4_11                              (cast_ready_pe_2_nw[4][11]),
    .merge_data_o_4_11                              (merge_data_nw_2_pe[4][11]),
    .merge_valid_o_4_11                             (merge_valid_nw_2_pe[4][11]),
    .merge_ready_i_4_11                             (merge_ready_pe_2_nw[4][11]),
    .gather_data_o_4_11                             (gather_data_nw_2_pe[4][11]),
    .gather_valid_o_4_11                            (gather_valid_nw_2_pe[4][11]),
    .gather_ready_i_4_11                            (gather_ready_pe_2_nw[4][11]),
    .cast_data_i_4_12                               (cast_data_pe_2_nw[4][12]),
    .cast_valid_i_4_12                              (cast_valid_pe_2_nw[4][12]),
    .cast_ready_o_4_12                              (cast_ready_nw_2_pe[4][12]),
    .merge_data_i_4_12                              (merge_data_pe_2_nw[4][12]),
    .merge_valid_i_4_12                             (merge_valid_pe_2_nw[4][12]),
    .merge_ready_o_4_12                             (merge_ready_nw_2_pe[4][12]),
    .gather_data_i_4_12                             (gather_data_pe_2_nw[4][12]),
    .gather_valid_i_4_12                            (gather_valid_pe_2_nw[4][12]),
    .gather_ready_o_4_12                            (gather_ready_nw_2_pe[4][12]),

    .cast_data_o_4_12                               (cast_data_nw_2_pe[4][12]),
    .cast_valid_o_4_12                              (cast_valid_nw_2_pe[4][12]),
    .cast_ready_i_4_12                              (cast_ready_pe_2_nw[4][12]),
    .merge_data_o_4_12                              (merge_data_nw_2_pe[4][12]),
    .merge_valid_o_4_12                             (merge_valid_nw_2_pe[4][12]),
    .merge_ready_i_4_12                             (merge_ready_pe_2_nw[4][12]),
    .gather_data_o_4_12                             (gather_data_nw_2_pe[4][12]),
    .gather_valid_o_4_12                            (gather_valid_nw_2_pe[4][12]),
    .gather_ready_i_4_12                            (gather_ready_pe_2_nw[4][12]),
    .cast_data_i_4_13                               (cast_data_pe_2_nw[4][13]),
    .cast_valid_i_4_13                              (cast_valid_pe_2_nw[4][13]),
    .cast_ready_o_4_13                              (cast_ready_nw_2_pe[4][13]),
    .merge_data_i_4_13                              (merge_data_pe_2_nw[4][13]),
    .merge_valid_i_4_13                             (merge_valid_pe_2_nw[4][13]),
    .merge_ready_o_4_13                             (merge_ready_nw_2_pe[4][13]),
    .gather_data_i_4_13                             (gather_data_pe_2_nw[4][13]),
    .gather_valid_i_4_13                            (gather_valid_pe_2_nw[4][13]),
    .gather_ready_o_4_13                            (gather_ready_nw_2_pe[4][13]),

    .cast_data_o_4_13                               (cast_data_nw_2_pe[4][13]),
    .cast_valid_o_4_13                              (cast_valid_nw_2_pe[4][13]),
    .cast_ready_i_4_13                              (cast_ready_pe_2_nw[4][13]),
    .merge_data_o_4_13                              (merge_data_nw_2_pe[4][13]),
    .merge_valid_o_4_13                             (merge_valid_nw_2_pe[4][13]),
    .merge_ready_i_4_13                             (merge_ready_pe_2_nw[4][13]),
    .gather_data_o_4_13                             (gather_data_nw_2_pe[4][13]),
    .gather_valid_o_4_13                            (gather_valid_nw_2_pe[4][13]),
    .gather_ready_i_4_13                            (gather_ready_pe_2_nw[4][13]),
    .cast_data_i_4_14                               (cast_data_pe_2_nw[4][14]),
    .cast_valid_i_4_14                              (cast_valid_pe_2_nw[4][14]),
    .cast_ready_o_4_14                              (cast_ready_nw_2_pe[4][14]),
    .merge_data_i_4_14                              (merge_data_pe_2_nw[4][14]),
    .merge_valid_i_4_14                             (merge_valid_pe_2_nw[4][14]),
    .merge_ready_o_4_14                             (merge_ready_nw_2_pe[4][14]),
    .gather_data_i_4_14                             (gather_data_pe_2_nw[4][14]),
    .gather_valid_i_4_14                            (gather_valid_pe_2_nw[4][14]),
    .gather_ready_o_4_14                            (gather_ready_nw_2_pe[4][14]),

    .cast_data_o_4_14                               (cast_data_nw_2_pe[4][14]),
    .cast_valid_o_4_14                              (cast_valid_nw_2_pe[4][14]),
    .cast_ready_i_4_14                              (cast_ready_pe_2_nw[4][14]),
    .merge_data_o_4_14                              (merge_data_nw_2_pe[4][14]),
    .merge_valid_o_4_14                             (merge_valid_nw_2_pe[4][14]),
    .merge_ready_i_4_14                             (merge_ready_pe_2_nw[4][14]),
    .gather_data_o_4_14                             (gather_data_nw_2_pe[4][14]),
    .gather_valid_o_4_14                            (gather_valid_nw_2_pe[4][14]),
    .gather_ready_i_4_14                            (gather_ready_pe_2_nw[4][14]),
    .cast_data_i_4_15                               (cast_data_pe_2_nw[4][15]),
    .cast_valid_i_4_15                              (cast_valid_pe_2_nw[4][15]),
    .cast_ready_o_4_15                              (cast_ready_nw_2_pe[4][15]),
    .merge_data_i_4_15                              (merge_data_pe_2_nw[4][15]),
    .merge_valid_i_4_15                             (merge_valid_pe_2_nw[4][15]),
    .merge_ready_o_4_15                             (merge_ready_nw_2_pe[4][15]),
    .gather_data_i_4_15                             (gather_data_pe_2_nw[4][15]),
    .gather_valid_i_4_15                            (gather_valid_pe_2_nw[4][15]),
    .gather_ready_o_4_15                            (gather_ready_nw_2_pe[4][15]),

    .cast_data_o_4_15                               (cast_data_nw_2_pe[4][15]),
    .cast_valid_o_4_15                              (cast_valid_nw_2_pe[4][15]),
    .cast_ready_i_4_15                              (cast_ready_pe_2_nw[4][15]),
    .merge_data_o_4_15                              (merge_data_nw_2_pe[4][15]),
    .merge_valid_o_4_15                             (merge_valid_nw_2_pe[4][15]),
    .merge_ready_i_4_15                             (merge_ready_pe_2_nw[4][15]),
    .gather_data_o_4_15                             (gather_data_nw_2_pe[4][15]),
    .gather_valid_o_4_15                            (gather_valid_nw_2_pe[4][15]),
    .gather_ready_i_4_15                            (gather_ready_pe_2_nw[4][15]),
    .cast_data_i_4_16                               (cast_data_pe_2_nw[4][16]),
    .cast_valid_i_4_16                              (cast_valid_pe_2_nw[4][16]),
    .cast_ready_o_4_16                              (cast_ready_nw_2_pe[4][16]),
    .merge_data_i_4_16                              (merge_data_pe_2_nw[4][16]),
    .merge_valid_i_4_16                             (merge_valid_pe_2_nw[4][16]),
    .merge_ready_o_4_16                             (merge_ready_nw_2_pe[4][16]),
    .gather_data_i_4_16                             (gather_data_pe_2_nw[4][16]),
    .gather_valid_i_4_16                            (gather_valid_pe_2_nw[4][16]),
    .gather_ready_o_4_16                            (gather_ready_nw_2_pe[4][16]),

    .cast_data_o_4_16                               (cast_data_nw_2_pe[4][16]),
    .cast_valid_o_4_16                              (cast_valid_nw_2_pe[4][16]),
    .cast_ready_i_4_16                              (cast_ready_pe_2_nw[4][16]),
    .merge_data_o_4_16                              (merge_data_nw_2_pe[4][16]),
    .merge_valid_o_4_16                             (merge_valid_nw_2_pe[4][16]),
    .merge_ready_i_4_16                             (merge_ready_pe_2_nw[4][16]),
    .gather_data_o_4_16                             (gather_data_nw_2_pe[4][16]),
    .gather_valid_o_4_16                            (gather_valid_nw_2_pe[4][16]),
    .gather_ready_i_4_16                            (gather_ready_pe_2_nw[4][16]),
    .cast_data_i_4_17                               (cast_data_pe_2_nw[4][17]),
    .cast_valid_i_4_17                              (cast_valid_pe_2_nw[4][17]),
    .cast_ready_o_4_17                              (cast_ready_nw_2_pe[4][17]),
    .merge_data_i_4_17                              (merge_data_pe_2_nw[4][17]),
    .merge_valid_i_4_17                             (merge_valid_pe_2_nw[4][17]),
    .merge_ready_o_4_17                             (merge_ready_nw_2_pe[4][17]),
    .gather_data_i_4_17                             (gather_data_pe_2_nw[4][17]),
    .gather_valid_i_4_17                            (gather_valid_pe_2_nw[4][17]),
    .gather_ready_o_4_17                            (gather_ready_nw_2_pe[4][17]),

    .cast_data_o_4_17                               (cast_data_nw_2_pe[4][17]),
    .cast_valid_o_4_17                              (cast_valid_nw_2_pe[4][17]),
    .cast_ready_i_4_17                              (cast_ready_pe_2_nw[4][17]),
    .merge_data_o_4_17                              (merge_data_nw_2_pe[4][17]),
    .merge_valid_o_4_17                             (merge_valid_nw_2_pe[4][17]),
    .merge_ready_i_4_17                             (merge_ready_pe_2_nw[4][17]),
    .gather_data_o_4_17                             (gather_data_nw_2_pe[4][17]),
    .gather_valid_o_4_17                            (gather_valid_nw_2_pe[4][17]),
    .gather_ready_i_4_17                            (gather_ready_pe_2_nw[4][17]),
    .cast_data_i_4_18                               (cast_data_pe_2_nw[4][18]),
    .cast_valid_i_4_18                              (cast_valid_pe_2_nw[4][18]),
    .cast_ready_o_4_18                              (cast_ready_nw_2_pe[4][18]),
    .merge_data_i_4_18                              (merge_data_pe_2_nw[4][18]),
    .merge_valid_i_4_18                             (merge_valid_pe_2_nw[4][18]),
    .merge_ready_o_4_18                             (merge_ready_nw_2_pe[4][18]),
    .gather_data_i_4_18                             (gather_data_pe_2_nw[4][18]),
    .gather_valid_i_4_18                            (gather_valid_pe_2_nw[4][18]),
    .gather_ready_o_4_18                            (gather_ready_nw_2_pe[4][18]),

    .cast_data_o_4_18                               (cast_data_nw_2_pe[4][18]),
    .cast_valid_o_4_18                              (cast_valid_nw_2_pe[4][18]),
    .cast_ready_i_4_18                              (cast_ready_pe_2_nw[4][18]),
    .merge_data_o_4_18                              (merge_data_nw_2_pe[4][18]),
    .merge_valid_o_4_18                             (merge_valid_nw_2_pe[4][18]),
    .merge_ready_i_4_18                             (merge_ready_pe_2_nw[4][18]),
    .gather_data_o_4_18                             (gather_data_nw_2_pe[4][18]),
    .gather_valid_o_4_18                            (gather_valid_nw_2_pe[4][18]),
    .gather_ready_i_4_18                            (gather_ready_pe_2_nw[4][18]),
    .cast_data_i_4_19                               (cast_data_pe_2_nw[4][19]),
    .cast_valid_i_4_19                              (cast_valid_pe_2_nw[4][19]),
    .cast_ready_o_4_19                              (cast_ready_nw_2_pe[4][19]),
    .merge_data_i_4_19                              (merge_data_pe_2_nw[4][19]),
    .merge_valid_i_4_19                             (merge_valid_pe_2_nw[4][19]),
    .merge_ready_o_4_19                             (merge_ready_nw_2_pe[4][19]),
    .gather_data_i_4_19                             (gather_data_pe_2_nw[4][19]),
    .gather_valid_i_4_19                            (gather_valid_pe_2_nw[4][19]),
    .gather_ready_o_4_19                            (gather_ready_nw_2_pe[4][19]),

    .cast_data_o_4_19                               (cast_data_nw_2_pe[4][19]),
    .cast_valid_o_4_19                              (cast_valid_nw_2_pe[4][19]),
    .cast_ready_i_4_19                              (cast_ready_pe_2_nw[4][19]),
    .merge_data_o_4_19                              (merge_data_nw_2_pe[4][19]),
    .merge_valid_o_4_19                             (merge_valid_nw_2_pe[4][19]),
    .merge_ready_i_4_19                             (merge_ready_pe_2_nw[4][19]),
    .gather_data_o_4_19                             (gather_data_nw_2_pe[4][19]),
    .gather_valid_o_4_19                            (gather_valid_nw_2_pe[4][19]),
    .gather_ready_i_4_19                            (gather_ready_pe_2_nw[4][19]),
    .cast_data_i_4_20                               (cast_data_pe_2_nw[4][20]),
    .cast_valid_i_4_20                              (cast_valid_pe_2_nw[4][20]),
    .cast_ready_o_4_20                              (cast_ready_nw_2_pe[4][20]),
    .merge_data_i_4_20                              (merge_data_pe_2_nw[4][20]),
    .merge_valid_i_4_20                             (merge_valid_pe_2_nw[4][20]),
    .merge_ready_o_4_20                             (merge_ready_nw_2_pe[4][20]),
    .gather_data_i_4_20                             (gather_data_pe_2_nw[4][20]),
    .gather_valid_i_4_20                            (gather_valid_pe_2_nw[4][20]),
    .gather_ready_o_4_20                            (gather_ready_nw_2_pe[4][20]),

    .cast_data_o_4_20                               (cast_data_nw_2_pe[4][20]),
    .cast_valid_o_4_20                              (cast_valid_nw_2_pe[4][20]),
    .cast_ready_i_4_20                              (cast_ready_pe_2_nw[4][20]),
    .merge_data_o_4_20                              (merge_data_nw_2_pe[4][20]),
    .merge_valid_o_4_20                             (merge_valid_nw_2_pe[4][20]),
    .merge_ready_i_4_20                             (merge_ready_pe_2_nw[4][20]),
    .gather_data_o_4_20                             (gather_data_nw_2_pe[4][20]),
    .gather_valid_o_4_20                            (gather_valid_nw_2_pe[4][20]),
    .gather_ready_i_4_20                            (gather_ready_pe_2_nw[4][20]),
    .cast_data_i_4_21                               (cast_data_pe_2_nw[4][21]),
    .cast_valid_i_4_21                              (cast_valid_pe_2_nw[4][21]),
    .cast_ready_o_4_21                              (cast_ready_nw_2_pe[4][21]),
    .merge_data_i_4_21                              (merge_data_pe_2_nw[4][21]),
    .merge_valid_i_4_21                             (merge_valid_pe_2_nw[4][21]),
    .merge_ready_o_4_21                             (merge_ready_nw_2_pe[4][21]),
    .gather_data_i_4_21                             (gather_data_pe_2_nw[4][21]),
    .gather_valid_i_4_21                            (gather_valid_pe_2_nw[4][21]),
    .gather_ready_o_4_21                            (gather_ready_nw_2_pe[4][21]),

    .cast_data_o_4_21                               (cast_data_nw_2_pe[4][21]),
    .cast_valid_o_4_21                              (cast_valid_nw_2_pe[4][21]),
    .cast_ready_i_4_21                              (cast_ready_pe_2_nw[4][21]),
    .merge_data_o_4_21                              (merge_data_nw_2_pe[4][21]),
    .merge_valid_o_4_21                             (merge_valid_nw_2_pe[4][21]),
    .merge_ready_i_4_21                             (merge_ready_pe_2_nw[4][21]),
    .gather_data_o_4_21                             (gather_data_nw_2_pe[4][21]),
    .gather_valid_o_4_21                            (gather_valid_nw_2_pe[4][21]),
    .gather_ready_i_4_21                            (gather_ready_pe_2_nw[4][21]),
    .cast_data_i_4_22                               (cast_data_pe_2_nw[4][22]),
    .cast_valid_i_4_22                              (cast_valid_pe_2_nw[4][22]),
    .cast_ready_o_4_22                              (cast_ready_nw_2_pe[4][22]),
    .merge_data_i_4_22                              (merge_data_pe_2_nw[4][22]),
    .merge_valid_i_4_22                             (merge_valid_pe_2_nw[4][22]),
    .merge_ready_o_4_22                             (merge_ready_nw_2_pe[4][22]),
    .gather_data_i_4_22                             (gather_data_pe_2_nw[4][22]),
    .gather_valid_i_4_22                            (gather_valid_pe_2_nw[4][22]),
    .gather_ready_o_4_22                            (gather_ready_nw_2_pe[4][22]),

    .cast_data_o_4_22                               (cast_data_nw_2_pe[4][22]),
    .cast_valid_o_4_22                              (cast_valid_nw_2_pe[4][22]),
    .cast_ready_i_4_22                              (cast_ready_pe_2_nw[4][22]),
    .merge_data_o_4_22                              (merge_data_nw_2_pe[4][22]),
    .merge_valid_o_4_22                             (merge_valid_nw_2_pe[4][22]),
    .merge_ready_i_4_22                             (merge_ready_pe_2_nw[4][22]),
    .gather_data_o_4_22                             (gather_data_nw_2_pe[4][22]),
    .gather_valid_o_4_22                            (gather_valid_nw_2_pe[4][22]),
    .gather_ready_i_4_22                            (gather_ready_pe_2_nw[4][22]),
    .cast_data_i_4_23                               (cast_data_pe_2_nw[4][23]),
    .cast_valid_i_4_23                              (cast_valid_pe_2_nw[4][23]),
    .cast_ready_o_4_23                              (cast_ready_nw_2_pe[4][23]),
    .merge_data_i_4_23                              (merge_data_pe_2_nw[4][23]),
    .merge_valid_i_4_23                             (merge_valid_pe_2_nw[4][23]),
    .merge_ready_o_4_23                             (merge_ready_nw_2_pe[4][23]),
    .gather_data_i_4_23                             (gather_data_pe_2_nw[4][23]),
    .gather_valid_i_4_23                            (gather_valid_pe_2_nw[4][23]),
    .gather_ready_o_4_23                            (gather_ready_nw_2_pe[4][23]),

    .cast_data_o_4_23                               (cast_data_nw_2_pe[4][23]),
    .cast_valid_o_4_23                              (cast_valid_nw_2_pe[4][23]),
    .cast_ready_i_4_23                              (cast_ready_pe_2_nw[4][23]),
    .merge_data_o_4_23                              (merge_data_nw_2_pe[4][23]),
    .merge_valid_o_4_23                             (merge_valid_nw_2_pe[4][23]),
    .merge_ready_i_4_23                             (merge_ready_pe_2_nw[4][23]),
    .gather_data_o_4_23                             (gather_data_nw_2_pe[4][23]),
    .gather_valid_o_4_23                            (gather_valid_nw_2_pe[4][23]),
    .gather_ready_i_4_23                            (gather_ready_pe_2_nw[4][23]),
    .cast_data_i_4_24                               (cast_data_pe_2_nw[4][24]),
    .cast_valid_i_4_24                              (cast_valid_pe_2_nw[4][24]),
    .cast_ready_o_4_24                              (cast_ready_nw_2_pe[4][24]),
    .merge_data_i_4_24                              (merge_data_pe_2_nw[4][24]),
    .merge_valid_i_4_24                             (merge_valid_pe_2_nw[4][24]),
    .merge_ready_o_4_24                             (merge_ready_nw_2_pe[4][24]),
    .gather_data_i_4_24                             (gather_data_pe_2_nw[4][24]),
    .gather_valid_i_4_24                            (gather_valid_pe_2_nw[4][24]),
    .gather_ready_o_4_24                            (gather_ready_nw_2_pe[4][24]),

    .cast_data_o_4_24                               (cast_data_nw_2_pe[4][24]),
    .cast_valid_o_4_24                              (cast_valid_nw_2_pe[4][24]),
    .cast_ready_i_4_24                              (cast_ready_pe_2_nw[4][24]),
    .merge_data_o_4_24                              (merge_data_nw_2_pe[4][24]),
    .merge_valid_o_4_24                             (merge_valid_nw_2_pe[4][24]),
    .merge_ready_i_4_24                             (merge_ready_pe_2_nw[4][24]),
    .gather_data_o_4_24                             (gather_data_nw_2_pe[4][24]),
    .gather_valid_o_4_24                            (gather_valid_nw_2_pe[4][24]),
    .gather_ready_i_4_24                            (gather_ready_pe_2_nw[4][24]),
    .cast_data_i_5_0                               (cast_data_pe_2_nw[5][0]),
    .cast_valid_i_5_0                              (cast_valid_pe_2_nw[5][0]),
    .cast_ready_o_5_0                              (cast_ready_nw_2_pe[5][0]),
    .merge_data_i_5_0                              (merge_data_pe_2_nw[5][0]),
    .merge_valid_i_5_0                             (merge_valid_pe_2_nw[5][0]),
    .merge_ready_o_5_0                             (merge_ready_nw_2_pe[5][0]),
    .gather_data_i_5_0                             (gather_data_pe_2_nw[5][0]),
    .gather_valid_i_5_0                            (gather_valid_pe_2_nw[5][0]),
    .gather_ready_o_5_0                            (gather_ready_nw_2_pe[5][0]),

    .cast_data_o_5_0                               (cast_data_nw_2_pe[5][0]),
    .cast_valid_o_5_0                              (cast_valid_nw_2_pe[5][0]),
    .cast_ready_i_5_0                              (cast_ready_pe_2_nw[5][0]),
    .merge_data_o_5_0                              (merge_data_nw_2_pe[5][0]),
    .merge_valid_o_5_0                             (merge_valid_nw_2_pe[5][0]),
    .merge_ready_i_5_0                             (merge_ready_pe_2_nw[5][0]),
    .gather_data_o_5_0                             (gather_data_nw_2_pe[5][0]),
    .gather_valid_o_5_0                            (gather_valid_nw_2_pe[5][0]),
    .gather_ready_i_5_0                            (gather_ready_pe_2_nw[5][0]),
    .cast_data_i_5_1                               (cast_data_pe_2_nw[5][1]),
    .cast_valid_i_5_1                              (cast_valid_pe_2_nw[5][1]),
    .cast_ready_o_5_1                              (cast_ready_nw_2_pe[5][1]),
    .merge_data_i_5_1                              (merge_data_pe_2_nw[5][1]),
    .merge_valid_i_5_1                             (merge_valid_pe_2_nw[5][1]),
    .merge_ready_o_5_1                             (merge_ready_nw_2_pe[5][1]),
    .gather_data_i_5_1                             (gather_data_pe_2_nw[5][1]),
    .gather_valid_i_5_1                            (gather_valid_pe_2_nw[5][1]),
    .gather_ready_o_5_1                            (gather_ready_nw_2_pe[5][1]),

    .cast_data_o_5_1                               (cast_data_nw_2_pe[5][1]),
    .cast_valid_o_5_1                              (cast_valid_nw_2_pe[5][1]),
    .cast_ready_i_5_1                              (cast_ready_pe_2_nw[5][1]),
    .merge_data_o_5_1                              (merge_data_nw_2_pe[5][1]),
    .merge_valid_o_5_1                             (merge_valid_nw_2_pe[5][1]),
    .merge_ready_i_5_1                             (merge_ready_pe_2_nw[5][1]),
    .gather_data_o_5_1                             (gather_data_nw_2_pe[5][1]),
    .gather_valid_o_5_1                            (gather_valid_nw_2_pe[5][1]),
    .gather_ready_i_5_1                            (gather_ready_pe_2_nw[5][1]),
    .cast_data_i_5_2                               (cast_data_pe_2_nw[5][2]),
    .cast_valid_i_5_2                              (cast_valid_pe_2_nw[5][2]),
    .cast_ready_o_5_2                              (cast_ready_nw_2_pe[5][2]),
    .merge_data_i_5_2                              (merge_data_pe_2_nw[5][2]),
    .merge_valid_i_5_2                             (merge_valid_pe_2_nw[5][2]),
    .merge_ready_o_5_2                             (merge_ready_nw_2_pe[5][2]),
    .gather_data_i_5_2                             (gather_data_pe_2_nw[5][2]),
    .gather_valid_i_5_2                            (gather_valid_pe_2_nw[5][2]),
    .gather_ready_o_5_2                            (gather_ready_nw_2_pe[5][2]),

    .cast_data_o_5_2                               (cast_data_nw_2_pe[5][2]),
    .cast_valid_o_5_2                              (cast_valid_nw_2_pe[5][2]),
    .cast_ready_i_5_2                              (cast_ready_pe_2_nw[5][2]),
    .merge_data_o_5_2                              (merge_data_nw_2_pe[5][2]),
    .merge_valid_o_5_2                             (merge_valid_nw_2_pe[5][2]),
    .merge_ready_i_5_2                             (merge_ready_pe_2_nw[5][2]),
    .gather_data_o_5_2                             (gather_data_nw_2_pe[5][2]),
    .gather_valid_o_5_2                            (gather_valid_nw_2_pe[5][2]),
    .gather_ready_i_5_2                            (gather_ready_pe_2_nw[5][2]),
    .cast_data_i_5_3                               (cast_data_pe_2_nw[5][3]),
    .cast_valid_i_5_3                              (cast_valid_pe_2_nw[5][3]),
    .cast_ready_o_5_3                              (cast_ready_nw_2_pe[5][3]),
    .merge_data_i_5_3                              (merge_data_pe_2_nw[5][3]),
    .merge_valid_i_5_3                             (merge_valid_pe_2_nw[5][3]),
    .merge_ready_o_5_3                             (merge_ready_nw_2_pe[5][3]),
    .gather_data_i_5_3                             (gather_data_pe_2_nw[5][3]),
    .gather_valid_i_5_3                            (gather_valid_pe_2_nw[5][3]),
    .gather_ready_o_5_3                            (gather_ready_nw_2_pe[5][3]),

    .cast_data_o_5_3                               (cast_data_nw_2_pe[5][3]),
    .cast_valid_o_5_3                              (cast_valid_nw_2_pe[5][3]),
    .cast_ready_i_5_3                              (cast_ready_pe_2_nw[5][3]),
    .merge_data_o_5_3                              (merge_data_nw_2_pe[5][3]),
    .merge_valid_o_5_3                             (merge_valid_nw_2_pe[5][3]),
    .merge_ready_i_5_3                             (merge_ready_pe_2_nw[5][3]),
    .gather_data_o_5_3                             (gather_data_nw_2_pe[5][3]),
    .gather_valid_o_5_3                            (gather_valid_nw_2_pe[5][3]),
    .gather_ready_i_5_3                            (gather_ready_pe_2_nw[5][3]),
    .cast_data_i_5_4                               (cast_data_pe_2_nw[5][4]),
    .cast_valid_i_5_4                              (cast_valid_pe_2_nw[5][4]),
    .cast_ready_o_5_4                              (cast_ready_nw_2_pe[5][4]),
    .merge_data_i_5_4                              (merge_data_pe_2_nw[5][4]),
    .merge_valid_i_5_4                             (merge_valid_pe_2_nw[5][4]),
    .merge_ready_o_5_4                             (merge_ready_nw_2_pe[5][4]),
    .gather_data_i_5_4                             (gather_data_pe_2_nw[5][4]),
    .gather_valid_i_5_4                            (gather_valid_pe_2_nw[5][4]),
    .gather_ready_o_5_4                            (gather_ready_nw_2_pe[5][4]),

    .cast_data_o_5_4                               (cast_data_nw_2_pe[5][4]),
    .cast_valid_o_5_4                              (cast_valid_nw_2_pe[5][4]),
    .cast_ready_i_5_4                              (cast_ready_pe_2_nw[5][4]),
    .merge_data_o_5_4                              (merge_data_nw_2_pe[5][4]),
    .merge_valid_o_5_4                             (merge_valid_nw_2_pe[5][4]),
    .merge_ready_i_5_4                             (merge_ready_pe_2_nw[5][4]),
    .gather_data_o_5_4                             (gather_data_nw_2_pe[5][4]),
    .gather_valid_o_5_4                            (gather_valid_nw_2_pe[5][4]),
    .gather_ready_i_5_4                            (gather_ready_pe_2_nw[5][4]),
    .cast_data_i_5_5                               (cast_data_pe_2_nw[5][5]),
    .cast_valid_i_5_5                              (cast_valid_pe_2_nw[5][5]),
    .cast_ready_o_5_5                              (cast_ready_nw_2_pe[5][5]),
    .merge_data_i_5_5                              (merge_data_pe_2_nw[5][5]),
    .merge_valid_i_5_5                             (merge_valid_pe_2_nw[5][5]),
    .merge_ready_o_5_5                             (merge_ready_nw_2_pe[5][5]),
    .gather_data_i_5_5                             (gather_data_pe_2_nw[5][5]),
    .gather_valid_i_5_5                            (gather_valid_pe_2_nw[5][5]),
    .gather_ready_o_5_5                            (gather_ready_nw_2_pe[5][5]),

    .cast_data_o_5_5                               (cast_data_nw_2_pe[5][5]),
    .cast_valid_o_5_5                              (cast_valid_nw_2_pe[5][5]),
    .cast_ready_i_5_5                              (cast_ready_pe_2_nw[5][5]),
    .merge_data_o_5_5                              (merge_data_nw_2_pe[5][5]),
    .merge_valid_o_5_5                             (merge_valid_nw_2_pe[5][5]),
    .merge_ready_i_5_5                             (merge_ready_pe_2_nw[5][5]),
    .gather_data_o_5_5                             (gather_data_nw_2_pe[5][5]),
    .gather_valid_o_5_5                            (gather_valid_nw_2_pe[5][5]),
    .gather_ready_i_5_5                            (gather_ready_pe_2_nw[5][5]),
    .cast_data_i_5_6                               (cast_data_pe_2_nw[5][6]),
    .cast_valid_i_5_6                              (cast_valid_pe_2_nw[5][6]),
    .cast_ready_o_5_6                              (cast_ready_nw_2_pe[5][6]),
    .merge_data_i_5_6                              (merge_data_pe_2_nw[5][6]),
    .merge_valid_i_5_6                             (merge_valid_pe_2_nw[5][6]),
    .merge_ready_o_5_6                             (merge_ready_nw_2_pe[5][6]),
    .gather_data_i_5_6                             (gather_data_pe_2_nw[5][6]),
    .gather_valid_i_5_6                            (gather_valid_pe_2_nw[5][6]),
    .gather_ready_o_5_6                            (gather_ready_nw_2_pe[5][6]),

    .cast_data_o_5_6                               (cast_data_nw_2_pe[5][6]),
    .cast_valid_o_5_6                              (cast_valid_nw_2_pe[5][6]),
    .cast_ready_i_5_6                              (cast_ready_pe_2_nw[5][6]),
    .merge_data_o_5_6                              (merge_data_nw_2_pe[5][6]),
    .merge_valid_o_5_6                             (merge_valid_nw_2_pe[5][6]),
    .merge_ready_i_5_6                             (merge_ready_pe_2_nw[5][6]),
    .gather_data_o_5_6                             (gather_data_nw_2_pe[5][6]),
    .gather_valid_o_5_6                            (gather_valid_nw_2_pe[5][6]),
    .gather_ready_i_5_6                            (gather_ready_pe_2_nw[5][6]),
    .cast_data_i_5_7                               (cast_data_pe_2_nw[5][7]),
    .cast_valid_i_5_7                              (cast_valid_pe_2_nw[5][7]),
    .cast_ready_o_5_7                              (cast_ready_nw_2_pe[5][7]),
    .merge_data_i_5_7                              (merge_data_pe_2_nw[5][7]),
    .merge_valid_i_5_7                             (merge_valid_pe_2_nw[5][7]),
    .merge_ready_o_5_7                             (merge_ready_nw_2_pe[5][7]),
    .gather_data_i_5_7                             (gather_data_pe_2_nw[5][7]),
    .gather_valid_i_5_7                            (gather_valid_pe_2_nw[5][7]),
    .gather_ready_o_5_7                            (gather_ready_nw_2_pe[5][7]),

    .cast_data_o_5_7                               (cast_data_nw_2_pe[5][7]),
    .cast_valid_o_5_7                              (cast_valid_nw_2_pe[5][7]),
    .cast_ready_i_5_7                              (cast_ready_pe_2_nw[5][7]),
    .merge_data_o_5_7                              (merge_data_nw_2_pe[5][7]),
    .merge_valid_o_5_7                             (merge_valid_nw_2_pe[5][7]),
    .merge_ready_i_5_7                             (merge_ready_pe_2_nw[5][7]),
    .gather_data_o_5_7                             (gather_data_nw_2_pe[5][7]),
    .gather_valid_o_5_7                            (gather_valid_nw_2_pe[5][7]),
    .gather_ready_i_5_7                            (gather_ready_pe_2_nw[5][7]),
    .cast_data_i_5_8                               (cast_data_pe_2_nw[5][8]),
    .cast_valid_i_5_8                              (cast_valid_pe_2_nw[5][8]),
    .cast_ready_o_5_8                              (cast_ready_nw_2_pe[5][8]),
    .merge_data_i_5_8                              (merge_data_pe_2_nw[5][8]),
    .merge_valid_i_5_8                             (merge_valid_pe_2_nw[5][8]),
    .merge_ready_o_5_8                             (merge_ready_nw_2_pe[5][8]),
    .gather_data_i_5_8                             (gather_data_pe_2_nw[5][8]),
    .gather_valid_i_5_8                            (gather_valid_pe_2_nw[5][8]),
    .gather_ready_o_5_8                            (gather_ready_nw_2_pe[5][8]),

    .cast_data_o_5_8                               (cast_data_nw_2_pe[5][8]),
    .cast_valid_o_5_8                              (cast_valid_nw_2_pe[5][8]),
    .cast_ready_i_5_8                              (cast_ready_pe_2_nw[5][8]),
    .merge_data_o_5_8                              (merge_data_nw_2_pe[5][8]),
    .merge_valid_o_5_8                             (merge_valid_nw_2_pe[5][8]),
    .merge_ready_i_5_8                             (merge_ready_pe_2_nw[5][8]),
    .gather_data_o_5_8                             (gather_data_nw_2_pe[5][8]),
    .gather_valid_o_5_8                            (gather_valid_nw_2_pe[5][8]),
    .gather_ready_i_5_8                            (gather_ready_pe_2_nw[5][8]),
    .cast_data_i_5_9                               (cast_data_pe_2_nw[5][9]),
    .cast_valid_i_5_9                              (cast_valid_pe_2_nw[5][9]),
    .cast_ready_o_5_9                              (cast_ready_nw_2_pe[5][9]),
    .merge_data_i_5_9                              (merge_data_pe_2_nw[5][9]),
    .merge_valid_i_5_9                             (merge_valid_pe_2_nw[5][9]),
    .merge_ready_o_5_9                             (merge_ready_nw_2_pe[5][9]),
    .gather_data_i_5_9                             (gather_data_pe_2_nw[5][9]),
    .gather_valid_i_5_9                            (gather_valid_pe_2_nw[5][9]),
    .gather_ready_o_5_9                            (gather_ready_nw_2_pe[5][9]),

    .cast_data_o_5_9                               (cast_data_nw_2_pe[5][9]),
    .cast_valid_o_5_9                              (cast_valid_nw_2_pe[5][9]),
    .cast_ready_i_5_9                              (cast_ready_pe_2_nw[5][9]),
    .merge_data_o_5_9                              (merge_data_nw_2_pe[5][9]),
    .merge_valid_o_5_9                             (merge_valid_nw_2_pe[5][9]),
    .merge_ready_i_5_9                             (merge_ready_pe_2_nw[5][9]),
    .gather_data_o_5_9                             (gather_data_nw_2_pe[5][9]),
    .gather_valid_o_5_9                            (gather_valid_nw_2_pe[5][9]),
    .gather_ready_i_5_9                            (gather_ready_pe_2_nw[5][9]),
    .cast_data_i_5_10                               (cast_data_pe_2_nw[5][10]),
    .cast_valid_i_5_10                              (cast_valid_pe_2_nw[5][10]),
    .cast_ready_o_5_10                              (cast_ready_nw_2_pe[5][10]),
    .merge_data_i_5_10                              (merge_data_pe_2_nw[5][10]),
    .merge_valid_i_5_10                             (merge_valid_pe_2_nw[5][10]),
    .merge_ready_o_5_10                             (merge_ready_nw_2_pe[5][10]),
    .gather_data_i_5_10                             (gather_data_pe_2_nw[5][10]),
    .gather_valid_i_5_10                            (gather_valid_pe_2_nw[5][10]),
    .gather_ready_o_5_10                            (gather_ready_nw_2_pe[5][10]),

    .cast_data_o_5_10                               (cast_data_nw_2_pe[5][10]),
    .cast_valid_o_5_10                              (cast_valid_nw_2_pe[5][10]),
    .cast_ready_i_5_10                              (cast_ready_pe_2_nw[5][10]),
    .merge_data_o_5_10                              (merge_data_nw_2_pe[5][10]),
    .merge_valid_o_5_10                             (merge_valid_nw_2_pe[5][10]),
    .merge_ready_i_5_10                             (merge_ready_pe_2_nw[5][10]),
    .gather_data_o_5_10                             (gather_data_nw_2_pe[5][10]),
    .gather_valid_o_5_10                            (gather_valid_nw_2_pe[5][10]),
    .gather_ready_i_5_10                            (gather_ready_pe_2_nw[5][10]),
    .cast_data_i_5_11                               (cast_data_pe_2_nw[5][11]),
    .cast_valid_i_5_11                              (cast_valid_pe_2_nw[5][11]),
    .cast_ready_o_5_11                              (cast_ready_nw_2_pe[5][11]),
    .merge_data_i_5_11                              (merge_data_pe_2_nw[5][11]),
    .merge_valid_i_5_11                             (merge_valid_pe_2_nw[5][11]),
    .merge_ready_o_5_11                             (merge_ready_nw_2_pe[5][11]),
    .gather_data_i_5_11                             (gather_data_pe_2_nw[5][11]),
    .gather_valid_i_5_11                            (gather_valid_pe_2_nw[5][11]),
    .gather_ready_o_5_11                            (gather_ready_nw_2_pe[5][11]),

    .cast_data_o_5_11                               (cast_data_nw_2_pe[5][11]),
    .cast_valid_o_5_11                              (cast_valid_nw_2_pe[5][11]),
    .cast_ready_i_5_11                              (cast_ready_pe_2_nw[5][11]),
    .merge_data_o_5_11                              (merge_data_nw_2_pe[5][11]),
    .merge_valid_o_5_11                             (merge_valid_nw_2_pe[5][11]),
    .merge_ready_i_5_11                             (merge_ready_pe_2_nw[5][11]),
    .gather_data_o_5_11                             (gather_data_nw_2_pe[5][11]),
    .gather_valid_o_5_11                            (gather_valid_nw_2_pe[5][11]),
    .gather_ready_i_5_11                            (gather_ready_pe_2_nw[5][11]),
    .cast_data_i_5_12                               (cast_data_pe_2_nw[5][12]),
    .cast_valid_i_5_12                              (cast_valid_pe_2_nw[5][12]),
    .cast_ready_o_5_12                              (cast_ready_nw_2_pe[5][12]),
    .merge_data_i_5_12                              (merge_data_pe_2_nw[5][12]),
    .merge_valid_i_5_12                             (merge_valid_pe_2_nw[5][12]),
    .merge_ready_o_5_12                             (merge_ready_nw_2_pe[5][12]),
    .gather_data_i_5_12                             (gather_data_pe_2_nw[5][12]),
    .gather_valid_i_5_12                            (gather_valid_pe_2_nw[5][12]),
    .gather_ready_o_5_12                            (gather_ready_nw_2_pe[5][12]),

    .cast_data_o_5_12                               (cast_data_nw_2_pe[5][12]),
    .cast_valid_o_5_12                              (cast_valid_nw_2_pe[5][12]),
    .cast_ready_i_5_12                              (cast_ready_pe_2_nw[5][12]),
    .merge_data_o_5_12                              (merge_data_nw_2_pe[5][12]),
    .merge_valid_o_5_12                             (merge_valid_nw_2_pe[5][12]),
    .merge_ready_i_5_12                             (merge_ready_pe_2_nw[5][12]),
    .gather_data_o_5_12                             (gather_data_nw_2_pe[5][12]),
    .gather_valid_o_5_12                            (gather_valid_nw_2_pe[5][12]),
    .gather_ready_i_5_12                            (gather_ready_pe_2_nw[5][12]),
    .cast_data_i_5_13                               (cast_data_pe_2_nw[5][13]),
    .cast_valid_i_5_13                              (cast_valid_pe_2_nw[5][13]),
    .cast_ready_o_5_13                              (cast_ready_nw_2_pe[5][13]),
    .merge_data_i_5_13                              (merge_data_pe_2_nw[5][13]),
    .merge_valid_i_5_13                             (merge_valid_pe_2_nw[5][13]),
    .merge_ready_o_5_13                             (merge_ready_nw_2_pe[5][13]),
    .gather_data_i_5_13                             (gather_data_pe_2_nw[5][13]),
    .gather_valid_i_5_13                            (gather_valid_pe_2_nw[5][13]),
    .gather_ready_o_5_13                            (gather_ready_nw_2_pe[5][13]),

    .cast_data_o_5_13                               (cast_data_nw_2_pe[5][13]),
    .cast_valid_o_5_13                              (cast_valid_nw_2_pe[5][13]),
    .cast_ready_i_5_13                              (cast_ready_pe_2_nw[5][13]),
    .merge_data_o_5_13                              (merge_data_nw_2_pe[5][13]),
    .merge_valid_o_5_13                             (merge_valid_nw_2_pe[5][13]),
    .merge_ready_i_5_13                             (merge_ready_pe_2_nw[5][13]),
    .gather_data_o_5_13                             (gather_data_nw_2_pe[5][13]),
    .gather_valid_o_5_13                            (gather_valid_nw_2_pe[5][13]),
    .gather_ready_i_5_13                            (gather_ready_pe_2_nw[5][13]),
    .cast_data_i_5_14                               (cast_data_pe_2_nw[5][14]),
    .cast_valid_i_5_14                              (cast_valid_pe_2_nw[5][14]),
    .cast_ready_o_5_14                              (cast_ready_nw_2_pe[5][14]),
    .merge_data_i_5_14                              (merge_data_pe_2_nw[5][14]),
    .merge_valid_i_5_14                             (merge_valid_pe_2_nw[5][14]),
    .merge_ready_o_5_14                             (merge_ready_nw_2_pe[5][14]),
    .gather_data_i_5_14                             (gather_data_pe_2_nw[5][14]),
    .gather_valid_i_5_14                            (gather_valid_pe_2_nw[5][14]),
    .gather_ready_o_5_14                            (gather_ready_nw_2_pe[5][14]),

    .cast_data_o_5_14                               (cast_data_nw_2_pe[5][14]),
    .cast_valid_o_5_14                              (cast_valid_nw_2_pe[5][14]),
    .cast_ready_i_5_14                              (cast_ready_pe_2_nw[5][14]),
    .merge_data_o_5_14                              (merge_data_nw_2_pe[5][14]),
    .merge_valid_o_5_14                             (merge_valid_nw_2_pe[5][14]),
    .merge_ready_i_5_14                             (merge_ready_pe_2_nw[5][14]),
    .gather_data_o_5_14                             (gather_data_nw_2_pe[5][14]),
    .gather_valid_o_5_14                            (gather_valid_nw_2_pe[5][14]),
    .gather_ready_i_5_14                            (gather_ready_pe_2_nw[5][14]),
    .cast_data_i_5_15                               (cast_data_pe_2_nw[5][15]),
    .cast_valid_i_5_15                              (cast_valid_pe_2_nw[5][15]),
    .cast_ready_o_5_15                              (cast_ready_nw_2_pe[5][15]),
    .merge_data_i_5_15                              (merge_data_pe_2_nw[5][15]),
    .merge_valid_i_5_15                             (merge_valid_pe_2_nw[5][15]),
    .merge_ready_o_5_15                             (merge_ready_nw_2_pe[5][15]),
    .gather_data_i_5_15                             (gather_data_pe_2_nw[5][15]),
    .gather_valid_i_5_15                            (gather_valid_pe_2_nw[5][15]),
    .gather_ready_o_5_15                            (gather_ready_nw_2_pe[5][15]),

    .cast_data_o_5_15                               (cast_data_nw_2_pe[5][15]),
    .cast_valid_o_5_15                              (cast_valid_nw_2_pe[5][15]),
    .cast_ready_i_5_15                              (cast_ready_pe_2_nw[5][15]),
    .merge_data_o_5_15                              (merge_data_nw_2_pe[5][15]),
    .merge_valid_o_5_15                             (merge_valid_nw_2_pe[5][15]),
    .merge_ready_i_5_15                             (merge_ready_pe_2_nw[5][15]),
    .gather_data_o_5_15                             (gather_data_nw_2_pe[5][15]),
    .gather_valid_o_5_15                            (gather_valid_nw_2_pe[5][15]),
    .gather_ready_i_5_15                            (gather_ready_pe_2_nw[5][15]),
    .cast_data_i_5_16                               (cast_data_pe_2_nw[5][16]),
    .cast_valid_i_5_16                              (cast_valid_pe_2_nw[5][16]),
    .cast_ready_o_5_16                              (cast_ready_nw_2_pe[5][16]),
    .merge_data_i_5_16                              (merge_data_pe_2_nw[5][16]),
    .merge_valid_i_5_16                             (merge_valid_pe_2_nw[5][16]),
    .merge_ready_o_5_16                             (merge_ready_nw_2_pe[5][16]),
    .gather_data_i_5_16                             (gather_data_pe_2_nw[5][16]),
    .gather_valid_i_5_16                            (gather_valid_pe_2_nw[5][16]),
    .gather_ready_o_5_16                            (gather_ready_nw_2_pe[5][16]),

    .cast_data_o_5_16                               (cast_data_nw_2_pe[5][16]),
    .cast_valid_o_5_16                              (cast_valid_nw_2_pe[5][16]),
    .cast_ready_i_5_16                              (cast_ready_pe_2_nw[5][16]),
    .merge_data_o_5_16                              (merge_data_nw_2_pe[5][16]),
    .merge_valid_o_5_16                             (merge_valid_nw_2_pe[5][16]),
    .merge_ready_i_5_16                             (merge_ready_pe_2_nw[5][16]),
    .gather_data_o_5_16                             (gather_data_nw_2_pe[5][16]),
    .gather_valid_o_5_16                            (gather_valid_nw_2_pe[5][16]),
    .gather_ready_i_5_16                            (gather_ready_pe_2_nw[5][16]),
    .cast_data_i_5_17                               (cast_data_pe_2_nw[5][17]),
    .cast_valid_i_5_17                              (cast_valid_pe_2_nw[5][17]),
    .cast_ready_o_5_17                              (cast_ready_nw_2_pe[5][17]),
    .merge_data_i_5_17                              (merge_data_pe_2_nw[5][17]),
    .merge_valid_i_5_17                             (merge_valid_pe_2_nw[5][17]),
    .merge_ready_o_5_17                             (merge_ready_nw_2_pe[5][17]),
    .gather_data_i_5_17                             (gather_data_pe_2_nw[5][17]),
    .gather_valid_i_5_17                            (gather_valid_pe_2_nw[5][17]),
    .gather_ready_o_5_17                            (gather_ready_nw_2_pe[5][17]),

    .cast_data_o_5_17                               (cast_data_nw_2_pe[5][17]),
    .cast_valid_o_5_17                              (cast_valid_nw_2_pe[5][17]),
    .cast_ready_i_5_17                              (cast_ready_pe_2_nw[5][17]),
    .merge_data_o_5_17                              (merge_data_nw_2_pe[5][17]),
    .merge_valid_o_5_17                             (merge_valid_nw_2_pe[5][17]),
    .merge_ready_i_5_17                             (merge_ready_pe_2_nw[5][17]),
    .gather_data_o_5_17                             (gather_data_nw_2_pe[5][17]),
    .gather_valid_o_5_17                            (gather_valid_nw_2_pe[5][17]),
    .gather_ready_i_5_17                            (gather_ready_pe_2_nw[5][17]),
    .cast_data_i_5_18                               (cast_data_pe_2_nw[5][18]),
    .cast_valid_i_5_18                              (cast_valid_pe_2_nw[5][18]),
    .cast_ready_o_5_18                              (cast_ready_nw_2_pe[5][18]),
    .merge_data_i_5_18                              (merge_data_pe_2_nw[5][18]),
    .merge_valid_i_5_18                             (merge_valid_pe_2_nw[5][18]),
    .merge_ready_o_5_18                             (merge_ready_nw_2_pe[5][18]),
    .gather_data_i_5_18                             (gather_data_pe_2_nw[5][18]),
    .gather_valid_i_5_18                            (gather_valid_pe_2_nw[5][18]),
    .gather_ready_o_5_18                            (gather_ready_nw_2_pe[5][18]),

    .cast_data_o_5_18                               (cast_data_nw_2_pe[5][18]),
    .cast_valid_o_5_18                              (cast_valid_nw_2_pe[5][18]),
    .cast_ready_i_5_18                              (cast_ready_pe_2_nw[5][18]),
    .merge_data_o_5_18                              (merge_data_nw_2_pe[5][18]),
    .merge_valid_o_5_18                             (merge_valid_nw_2_pe[5][18]),
    .merge_ready_i_5_18                             (merge_ready_pe_2_nw[5][18]),
    .gather_data_o_5_18                             (gather_data_nw_2_pe[5][18]),
    .gather_valid_o_5_18                            (gather_valid_nw_2_pe[5][18]),
    .gather_ready_i_5_18                            (gather_ready_pe_2_nw[5][18]),
    .cast_data_i_5_19                               (cast_data_pe_2_nw[5][19]),
    .cast_valid_i_5_19                              (cast_valid_pe_2_nw[5][19]),
    .cast_ready_o_5_19                              (cast_ready_nw_2_pe[5][19]),
    .merge_data_i_5_19                              (merge_data_pe_2_nw[5][19]),
    .merge_valid_i_5_19                             (merge_valid_pe_2_nw[5][19]),
    .merge_ready_o_5_19                             (merge_ready_nw_2_pe[5][19]),
    .gather_data_i_5_19                             (gather_data_pe_2_nw[5][19]),
    .gather_valid_i_5_19                            (gather_valid_pe_2_nw[5][19]),
    .gather_ready_o_5_19                            (gather_ready_nw_2_pe[5][19]),

    .cast_data_o_5_19                               (cast_data_nw_2_pe[5][19]),
    .cast_valid_o_5_19                              (cast_valid_nw_2_pe[5][19]),
    .cast_ready_i_5_19                              (cast_ready_pe_2_nw[5][19]),
    .merge_data_o_5_19                              (merge_data_nw_2_pe[5][19]),
    .merge_valid_o_5_19                             (merge_valid_nw_2_pe[5][19]),
    .merge_ready_i_5_19                             (merge_ready_pe_2_nw[5][19]),
    .gather_data_o_5_19                             (gather_data_nw_2_pe[5][19]),
    .gather_valid_o_5_19                            (gather_valid_nw_2_pe[5][19]),
    .gather_ready_i_5_19                            (gather_ready_pe_2_nw[5][19]),
    .cast_data_i_5_20                               (cast_data_pe_2_nw[5][20]),
    .cast_valid_i_5_20                              (cast_valid_pe_2_nw[5][20]),
    .cast_ready_o_5_20                              (cast_ready_nw_2_pe[5][20]),
    .merge_data_i_5_20                              (merge_data_pe_2_nw[5][20]),
    .merge_valid_i_5_20                             (merge_valid_pe_2_nw[5][20]),
    .merge_ready_o_5_20                             (merge_ready_nw_2_pe[5][20]),
    .gather_data_i_5_20                             (gather_data_pe_2_nw[5][20]),
    .gather_valid_i_5_20                            (gather_valid_pe_2_nw[5][20]),
    .gather_ready_o_5_20                            (gather_ready_nw_2_pe[5][20]),

    .cast_data_o_5_20                               (cast_data_nw_2_pe[5][20]),
    .cast_valid_o_5_20                              (cast_valid_nw_2_pe[5][20]),
    .cast_ready_i_5_20                              (cast_ready_pe_2_nw[5][20]),
    .merge_data_o_5_20                              (merge_data_nw_2_pe[5][20]),
    .merge_valid_o_5_20                             (merge_valid_nw_2_pe[5][20]),
    .merge_ready_i_5_20                             (merge_ready_pe_2_nw[5][20]),
    .gather_data_o_5_20                             (gather_data_nw_2_pe[5][20]),
    .gather_valid_o_5_20                            (gather_valid_nw_2_pe[5][20]),
    .gather_ready_i_5_20                            (gather_ready_pe_2_nw[5][20]),
    .cast_data_i_5_21                               (cast_data_pe_2_nw[5][21]),
    .cast_valid_i_5_21                              (cast_valid_pe_2_nw[5][21]),
    .cast_ready_o_5_21                              (cast_ready_nw_2_pe[5][21]),
    .merge_data_i_5_21                              (merge_data_pe_2_nw[5][21]),
    .merge_valid_i_5_21                             (merge_valid_pe_2_nw[5][21]),
    .merge_ready_o_5_21                             (merge_ready_nw_2_pe[5][21]),
    .gather_data_i_5_21                             (gather_data_pe_2_nw[5][21]),
    .gather_valid_i_5_21                            (gather_valid_pe_2_nw[5][21]),
    .gather_ready_o_5_21                            (gather_ready_nw_2_pe[5][21]),

    .cast_data_o_5_21                               (cast_data_nw_2_pe[5][21]),
    .cast_valid_o_5_21                              (cast_valid_nw_2_pe[5][21]),
    .cast_ready_i_5_21                              (cast_ready_pe_2_nw[5][21]),
    .merge_data_o_5_21                              (merge_data_nw_2_pe[5][21]),
    .merge_valid_o_5_21                             (merge_valid_nw_2_pe[5][21]),
    .merge_ready_i_5_21                             (merge_ready_pe_2_nw[5][21]),
    .gather_data_o_5_21                             (gather_data_nw_2_pe[5][21]),
    .gather_valid_o_5_21                            (gather_valid_nw_2_pe[5][21]),
    .gather_ready_i_5_21                            (gather_ready_pe_2_nw[5][21]),
    .cast_data_i_5_22                               (cast_data_pe_2_nw[5][22]),
    .cast_valid_i_5_22                              (cast_valid_pe_2_nw[5][22]),
    .cast_ready_o_5_22                              (cast_ready_nw_2_pe[5][22]),
    .merge_data_i_5_22                              (merge_data_pe_2_nw[5][22]),
    .merge_valid_i_5_22                             (merge_valid_pe_2_nw[5][22]),
    .merge_ready_o_5_22                             (merge_ready_nw_2_pe[5][22]),
    .gather_data_i_5_22                             (gather_data_pe_2_nw[5][22]),
    .gather_valid_i_5_22                            (gather_valid_pe_2_nw[5][22]),
    .gather_ready_o_5_22                            (gather_ready_nw_2_pe[5][22]),

    .cast_data_o_5_22                               (cast_data_nw_2_pe[5][22]),
    .cast_valid_o_5_22                              (cast_valid_nw_2_pe[5][22]),
    .cast_ready_i_5_22                              (cast_ready_pe_2_nw[5][22]),
    .merge_data_o_5_22                              (merge_data_nw_2_pe[5][22]),
    .merge_valid_o_5_22                             (merge_valid_nw_2_pe[5][22]),
    .merge_ready_i_5_22                             (merge_ready_pe_2_nw[5][22]),
    .gather_data_o_5_22                             (gather_data_nw_2_pe[5][22]),
    .gather_valid_o_5_22                            (gather_valid_nw_2_pe[5][22]),
    .gather_ready_i_5_22                            (gather_ready_pe_2_nw[5][22]),
    .cast_data_i_5_23                               (cast_data_pe_2_nw[5][23]),
    .cast_valid_i_5_23                              (cast_valid_pe_2_nw[5][23]),
    .cast_ready_o_5_23                              (cast_ready_nw_2_pe[5][23]),
    .merge_data_i_5_23                              (merge_data_pe_2_nw[5][23]),
    .merge_valid_i_5_23                             (merge_valid_pe_2_nw[5][23]),
    .merge_ready_o_5_23                             (merge_ready_nw_2_pe[5][23]),
    .gather_data_i_5_23                             (gather_data_pe_2_nw[5][23]),
    .gather_valid_i_5_23                            (gather_valid_pe_2_nw[5][23]),
    .gather_ready_o_5_23                            (gather_ready_nw_2_pe[5][23]),

    .cast_data_o_5_23                               (cast_data_nw_2_pe[5][23]),
    .cast_valid_o_5_23                              (cast_valid_nw_2_pe[5][23]),
    .cast_ready_i_5_23                              (cast_ready_pe_2_nw[5][23]),
    .merge_data_o_5_23                              (merge_data_nw_2_pe[5][23]),
    .merge_valid_o_5_23                             (merge_valid_nw_2_pe[5][23]),
    .merge_ready_i_5_23                             (merge_ready_pe_2_nw[5][23]),
    .gather_data_o_5_23                             (gather_data_nw_2_pe[5][23]),
    .gather_valid_o_5_23                            (gather_valid_nw_2_pe[5][23]),
    .gather_ready_i_5_23                            (gather_ready_pe_2_nw[5][23]),
    .cast_data_i_5_24                               (cast_data_pe_2_nw[5][24]),
    .cast_valid_i_5_24                              (cast_valid_pe_2_nw[5][24]),
    .cast_ready_o_5_24                              (cast_ready_nw_2_pe[5][24]),
    .merge_data_i_5_24                              (merge_data_pe_2_nw[5][24]),
    .merge_valid_i_5_24                             (merge_valid_pe_2_nw[5][24]),
    .merge_ready_o_5_24                             (merge_ready_nw_2_pe[5][24]),
    .gather_data_i_5_24                             (gather_data_pe_2_nw[5][24]),
    .gather_valid_i_5_24                            (gather_valid_pe_2_nw[5][24]),
    .gather_ready_o_5_24                            (gather_ready_nw_2_pe[5][24]),

    .cast_data_o_5_24                               (cast_data_nw_2_pe[5][24]),
    .cast_valid_o_5_24                              (cast_valid_nw_2_pe[5][24]),
    .cast_ready_i_5_24                              (cast_ready_pe_2_nw[5][24]),
    .merge_data_o_5_24                              (merge_data_nw_2_pe[5][24]),
    .merge_valid_o_5_24                             (merge_valid_nw_2_pe[5][24]),
    .merge_ready_i_5_24                             (merge_ready_pe_2_nw[5][24]),
    .gather_data_o_5_24                             (gather_data_nw_2_pe[5][24]),
    .gather_valid_o_5_24                            (gather_valid_nw_2_pe[5][24]),
    .gather_ready_i_5_24                            (gather_ready_pe_2_nw[5][24]),
    .cast_data_i_6_0                               (cast_data_pe_2_nw[6][0]),
    .cast_valid_i_6_0                              (cast_valid_pe_2_nw[6][0]),
    .cast_ready_o_6_0                              (cast_ready_nw_2_pe[6][0]),
    .merge_data_i_6_0                              (merge_data_pe_2_nw[6][0]),
    .merge_valid_i_6_0                             (merge_valid_pe_2_nw[6][0]),
    .merge_ready_o_6_0                             (merge_ready_nw_2_pe[6][0]),
    .gather_data_i_6_0                             (gather_data_pe_2_nw[6][0]),
    .gather_valid_i_6_0                            (gather_valid_pe_2_nw[6][0]),
    .gather_ready_o_6_0                            (gather_ready_nw_2_pe[6][0]),

    .cast_data_o_6_0                               (cast_data_nw_2_pe[6][0]),
    .cast_valid_o_6_0                              (cast_valid_nw_2_pe[6][0]),
    .cast_ready_i_6_0                              (cast_ready_pe_2_nw[6][0]),
    .merge_data_o_6_0                              (merge_data_nw_2_pe[6][0]),
    .merge_valid_o_6_0                             (merge_valid_nw_2_pe[6][0]),
    .merge_ready_i_6_0                             (merge_ready_pe_2_nw[6][0]),
    .gather_data_o_6_0                             (gather_data_nw_2_pe[6][0]),
    .gather_valid_o_6_0                            (gather_valid_nw_2_pe[6][0]),
    .gather_ready_i_6_0                            (gather_ready_pe_2_nw[6][0]),
    .cast_data_i_6_1                               (cast_data_pe_2_nw[6][1]),
    .cast_valid_i_6_1                              (cast_valid_pe_2_nw[6][1]),
    .cast_ready_o_6_1                              (cast_ready_nw_2_pe[6][1]),
    .merge_data_i_6_1                              (merge_data_pe_2_nw[6][1]),
    .merge_valid_i_6_1                             (merge_valid_pe_2_nw[6][1]),
    .merge_ready_o_6_1                             (merge_ready_nw_2_pe[6][1]),
    .gather_data_i_6_1                             (gather_data_pe_2_nw[6][1]),
    .gather_valid_i_6_1                            (gather_valid_pe_2_nw[6][1]),
    .gather_ready_o_6_1                            (gather_ready_nw_2_pe[6][1]),

    .cast_data_o_6_1                               (cast_data_nw_2_pe[6][1]),
    .cast_valid_o_6_1                              (cast_valid_nw_2_pe[6][1]),
    .cast_ready_i_6_1                              (cast_ready_pe_2_nw[6][1]),
    .merge_data_o_6_1                              (merge_data_nw_2_pe[6][1]),
    .merge_valid_o_6_1                             (merge_valid_nw_2_pe[6][1]),
    .merge_ready_i_6_1                             (merge_ready_pe_2_nw[6][1]),
    .gather_data_o_6_1                             (gather_data_nw_2_pe[6][1]),
    .gather_valid_o_6_1                            (gather_valid_nw_2_pe[6][1]),
    .gather_ready_i_6_1                            (gather_ready_pe_2_nw[6][1]),
    .cast_data_i_6_2                               (cast_data_pe_2_nw[6][2]),
    .cast_valid_i_6_2                              (cast_valid_pe_2_nw[6][2]),
    .cast_ready_o_6_2                              (cast_ready_nw_2_pe[6][2]),
    .merge_data_i_6_2                              (merge_data_pe_2_nw[6][2]),
    .merge_valid_i_6_2                             (merge_valid_pe_2_nw[6][2]),
    .merge_ready_o_6_2                             (merge_ready_nw_2_pe[6][2]),
    .gather_data_i_6_2                             (gather_data_pe_2_nw[6][2]),
    .gather_valid_i_6_2                            (gather_valid_pe_2_nw[6][2]),
    .gather_ready_o_6_2                            (gather_ready_nw_2_pe[6][2]),

    .cast_data_o_6_2                               (cast_data_nw_2_pe[6][2]),
    .cast_valid_o_6_2                              (cast_valid_nw_2_pe[6][2]),
    .cast_ready_i_6_2                              (cast_ready_pe_2_nw[6][2]),
    .merge_data_o_6_2                              (merge_data_nw_2_pe[6][2]),
    .merge_valid_o_6_2                             (merge_valid_nw_2_pe[6][2]),
    .merge_ready_i_6_2                             (merge_ready_pe_2_nw[6][2]),
    .gather_data_o_6_2                             (gather_data_nw_2_pe[6][2]),
    .gather_valid_o_6_2                            (gather_valid_nw_2_pe[6][2]),
    .gather_ready_i_6_2                            (gather_ready_pe_2_nw[6][2]),
    .cast_data_i_6_3                               (cast_data_pe_2_nw[6][3]),
    .cast_valid_i_6_3                              (cast_valid_pe_2_nw[6][3]),
    .cast_ready_o_6_3                              (cast_ready_nw_2_pe[6][3]),
    .merge_data_i_6_3                              (merge_data_pe_2_nw[6][3]),
    .merge_valid_i_6_3                             (merge_valid_pe_2_nw[6][3]),
    .merge_ready_o_6_3                             (merge_ready_nw_2_pe[6][3]),
    .gather_data_i_6_3                             (gather_data_pe_2_nw[6][3]),
    .gather_valid_i_6_3                            (gather_valid_pe_2_nw[6][3]),
    .gather_ready_o_6_3                            (gather_ready_nw_2_pe[6][3]),

    .cast_data_o_6_3                               (cast_data_nw_2_pe[6][3]),
    .cast_valid_o_6_3                              (cast_valid_nw_2_pe[6][3]),
    .cast_ready_i_6_3                              (cast_ready_pe_2_nw[6][3]),
    .merge_data_o_6_3                              (merge_data_nw_2_pe[6][3]),
    .merge_valid_o_6_3                             (merge_valid_nw_2_pe[6][3]),
    .merge_ready_i_6_3                             (merge_ready_pe_2_nw[6][3]),
    .gather_data_o_6_3                             (gather_data_nw_2_pe[6][3]),
    .gather_valid_o_6_3                            (gather_valid_nw_2_pe[6][3]),
    .gather_ready_i_6_3                            (gather_ready_pe_2_nw[6][3]),
    .cast_data_i_6_4                               (cast_data_pe_2_nw[6][4]),
    .cast_valid_i_6_4                              (cast_valid_pe_2_nw[6][4]),
    .cast_ready_o_6_4                              (cast_ready_nw_2_pe[6][4]),
    .merge_data_i_6_4                              (merge_data_pe_2_nw[6][4]),
    .merge_valid_i_6_4                             (merge_valid_pe_2_nw[6][4]),
    .merge_ready_o_6_4                             (merge_ready_nw_2_pe[6][4]),
    .gather_data_i_6_4                             (gather_data_pe_2_nw[6][4]),
    .gather_valid_i_6_4                            (gather_valid_pe_2_nw[6][4]),
    .gather_ready_o_6_4                            (gather_ready_nw_2_pe[6][4]),

    .cast_data_o_6_4                               (cast_data_nw_2_pe[6][4]),
    .cast_valid_o_6_4                              (cast_valid_nw_2_pe[6][4]),
    .cast_ready_i_6_4                              (cast_ready_pe_2_nw[6][4]),
    .merge_data_o_6_4                              (merge_data_nw_2_pe[6][4]),
    .merge_valid_o_6_4                             (merge_valid_nw_2_pe[6][4]),
    .merge_ready_i_6_4                             (merge_ready_pe_2_nw[6][4]),
    .gather_data_o_6_4                             (gather_data_nw_2_pe[6][4]),
    .gather_valid_o_6_4                            (gather_valid_nw_2_pe[6][4]),
    .gather_ready_i_6_4                            (gather_ready_pe_2_nw[6][4]),
    .cast_data_i_6_5                               (cast_data_pe_2_nw[6][5]),
    .cast_valid_i_6_5                              (cast_valid_pe_2_nw[6][5]),
    .cast_ready_o_6_5                              (cast_ready_nw_2_pe[6][5]),
    .merge_data_i_6_5                              (merge_data_pe_2_nw[6][5]),
    .merge_valid_i_6_5                             (merge_valid_pe_2_nw[6][5]),
    .merge_ready_o_6_5                             (merge_ready_nw_2_pe[6][5]),
    .gather_data_i_6_5                             (gather_data_pe_2_nw[6][5]),
    .gather_valid_i_6_5                            (gather_valid_pe_2_nw[6][5]),
    .gather_ready_o_6_5                            (gather_ready_nw_2_pe[6][5]),

    .cast_data_o_6_5                               (cast_data_nw_2_pe[6][5]),
    .cast_valid_o_6_5                              (cast_valid_nw_2_pe[6][5]),
    .cast_ready_i_6_5                              (cast_ready_pe_2_nw[6][5]),
    .merge_data_o_6_5                              (merge_data_nw_2_pe[6][5]),
    .merge_valid_o_6_5                             (merge_valid_nw_2_pe[6][5]),
    .merge_ready_i_6_5                             (merge_ready_pe_2_nw[6][5]),
    .gather_data_o_6_5                             (gather_data_nw_2_pe[6][5]),
    .gather_valid_o_6_5                            (gather_valid_nw_2_pe[6][5]),
    .gather_ready_i_6_5                            (gather_ready_pe_2_nw[6][5]),
    .cast_data_i_6_6                               (cast_data_pe_2_nw[6][6]),
    .cast_valid_i_6_6                              (cast_valid_pe_2_nw[6][6]),
    .cast_ready_o_6_6                              (cast_ready_nw_2_pe[6][6]),
    .merge_data_i_6_6                              (merge_data_pe_2_nw[6][6]),
    .merge_valid_i_6_6                             (merge_valid_pe_2_nw[6][6]),
    .merge_ready_o_6_6                             (merge_ready_nw_2_pe[6][6]),
    .gather_data_i_6_6                             (gather_data_pe_2_nw[6][6]),
    .gather_valid_i_6_6                            (gather_valid_pe_2_nw[6][6]),
    .gather_ready_o_6_6                            (gather_ready_nw_2_pe[6][6]),

    .cast_data_o_6_6                               (cast_data_nw_2_pe[6][6]),
    .cast_valid_o_6_6                              (cast_valid_nw_2_pe[6][6]),
    .cast_ready_i_6_6                              (cast_ready_pe_2_nw[6][6]),
    .merge_data_o_6_6                              (merge_data_nw_2_pe[6][6]),
    .merge_valid_o_6_6                             (merge_valid_nw_2_pe[6][6]),
    .merge_ready_i_6_6                             (merge_ready_pe_2_nw[6][6]),
    .gather_data_o_6_6                             (gather_data_nw_2_pe[6][6]),
    .gather_valid_o_6_6                            (gather_valid_nw_2_pe[6][6]),
    .gather_ready_i_6_6                            (gather_ready_pe_2_nw[6][6]),
    .cast_data_i_6_7                               (cast_data_pe_2_nw[6][7]),
    .cast_valid_i_6_7                              (cast_valid_pe_2_nw[6][7]),
    .cast_ready_o_6_7                              (cast_ready_nw_2_pe[6][7]),
    .merge_data_i_6_7                              (merge_data_pe_2_nw[6][7]),
    .merge_valid_i_6_7                             (merge_valid_pe_2_nw[6][7]),
    .merge_ready_o_6_7                             (merge_ready_nw_2_pe[6][7]),
    .gather_data_i_6_7                             (gather_data_pe_2_nw[6][7]),
    .gather_valid_i_6_7                            (gather_valid_pe_2_nw[6][7]),
    .gather_ready_o_6_7                            (gather_ready_nw_2_pe[6][7]),

    .cast_data_o_6_7                               (cast_data_nw_2_pe[6][7]),
    .cast_valid_o_6_7                              (cast_valid_nw_2_pe[6][7]),
    .cast_ready_i_6_7                              (cast_ready_pe_2_nw[6][7]),
    .merge_data_o_6_7                              (merge_data_nw_2_pe[6][7]),
    .merge_valid_o_6_7                             (merge_valid_nw_2_pe[6][7]),
    .merge_ready_i_6_7                             (merge_ready_pe_2_nw[6][7]),
    .gather_data_o_6_7                             (gather_data_nw_2_pe[6][7]),
    .gather_valid_o_6_7                            (gather_valid_nw_2_pe[6][7]),
    .gather_ready_i_6_7                            (gather_ready_pe_2_nw[6][7]),
    .cast_data_i_6_8                               (cast_data_pe_2_nw[6][8]),
    .cast_valid_i_6_8                              (cast_valid_pe_2_nw[6][8]),
    .cast_ready_o_6_8                              (cast_ready_nw_2_pe[6][8]),
    .merge_data_i_6_8                              (merge_data_pe_2_nw[6][8]),
    .merge_valid_i_6_8                             (merge_valid_pe_2_nw[6][8]),
    .merge_ready_o_6_8                             (merge_ready_nw_2_pe[6][8]),
    .gather_data_i_6_8                             (gather_data_pe_2_nw[6][8]),
    .gather_valid_i_6_8                            (gather_valid_pe_2_nw[6][8]),
    .gather_ready_o_6_8                            (gather_ready_nw_2_pe[6][8]),

    .cast_data_o_6_8                               (cast_data_nw_2_pe[6][8]),
    .cast_valid_o_6_8                              (cast_valid_nw_2_pe[6][8]),
    .cast_ready_i_6_8                              (cast_ready_pe_2_nw[6][8]),
    .merge_data_o_6_8                              (merge_data_nw_2_pe[6][8]),
    .merge_valid_o_6_8                             (merge_valid_nw_2_pe[6][8]),
    .merge_ready_i_6_8                             (merge_ready_pe_2_nw[6][8]),
    .gather_data_o_6_8                             (gather_data_nw_2_pe[6][8]),
    .gather_valid_o_6_8                            (gather_valid_nw_2_pe[6][8]),
    .gather_ready_i_6_8                            (gather_ready_pe_2_nw[6][8]),
    .cast_data_i_6_9                               (cast_data_pe_2_nw[6][9]),
    .cast_valid_i_6_9                              (cast_valid_pe_2_nw[6][9]),
    .cast_ready_o_6_9                              (cast_ready_nw_2_pe[6][9]),
    .merge_data_i_6_9                              (merge_data_pe_2_nw[6][9]),
    .merge_valid_i_6_9                             (merge_valid_pe_2_nw[6][9]),
    .merge_ready_o_6_9                             (merge_ready_nw_2_pe[6][9]),
    .gather_data_i_6_9                             (gather_data_pe_2_nw[6][9]),
    .gather_valid_i_6_9                            (gather_valid_pe_2_nw[6][9]),
    .gather_ready_o_6_9                            (gather_ready_nw_2_pe[6][9]),

    .cast_data_o_6_9                               (cast_data_nw_2_pe[6][9]),
    .cast_valid_o_6_9                              (cast_valid_nw_2_pe[6][9]),
    .cast_ready_i_6_9                              (cast_ready_pe_2_nw[6][9]),
    .merge_data_o_6_9                              (merge_data_nw_2_pe[6][9]),
    .merge_valid_o_6_9                             (merge_valid_nw_2_pe[6][9]),
    .merge_ready_i_6_9                             (merge_ready_pe_2_nw[6][9]),
    .gather_data_o_6_9                             (gather_data_nw_2_pe[6][9]),
    .gather_valid_o_6_9                            (gather_valid_nw_2_pe[6][9]),
    .gather_ready_i_6_9                            (gather_ready_pe_2_nw[6][9]),
    .cast_data_i_6_10                               (cast_data_pe_2_nw[6][10]),
    .cast_valid_i_6_10                              (cast_valid_pe_2_nw[6][10]),
    .cast_ready_o_6_10                              (cast_ready_nw_2_pe[6][10]),
    .merge_data_i_6_10                              (merge_data_pe_2_nw[6][10]),
    .merge_valid_i_6_10                             (merge_valid_pe_2_nw[6][10]),
    .merge_ready_o_6_10                             (merge_ready_nw_2_pe[6][10]),
    .gather_data_i_6_10                             (gather_data_pe_2_nw[6][10]),
    .gather_valid_i_6_10                            (gather_valid_pe_2_nw[6][10]),
    .gather_ready_o_6_10                            (gather_ready_nw_2_pe[6][10]),

    .cast_data_o_6_10                               (cast_data_nw_2_pe[6][10]),
    .cast_valid_o_6_10                              (cast_valid_nw_2_pe[6][10]),
    .cast_ready_i_6_10                              (cast_ready_pe_2_nw[6][10]),
    .merge_data_o_6_10                              (merge_data_nw_2_pe[6][10]),
    .merge_valid_o_6_10                             (merge_valid_nw_2_pe[6][10]),
    .merge_ready_i_6_10                             (merge_ready_pe_2_nw[6][10]),
    .gather_data_o_6_10                             (gather_data_nw_2_pe[6][10]),
    .gather_valid_o_6_10                            (gather_valid_nw_2_pe[6][10]),
    .gather_ready_i_6_10                            (gather_ready_pe_2_nw[6][10]),
    .cast_data_i_6_11                               (cast_data_pe_2_nw[6][11]),
    .cast_valid_i_6_11                              (cast_valid_pe_2_nw[6][11]),
    .cast_ready_o_6_11                              (cast_ready_nw_2_pe[6][11]),
    .merge_data_i_6_11                              (merge_data_pe_2_nw[6][11]),
    .merge_valid_i_6_11                             (merge_valid_pe_2_nw[6][11]),
    .merge_ready_o_6_11                             (merge_ready_nw_2_pe[6][11]),
    .gather_data_i_6_11                             (gather_data_pe_2_nw[6][11]),
    .gather_valid_i_6_11                            (gather_valid_pe_2_nw[6][11]),
    .gather_ready_o_6_11                            (gather_ready_nw_2_pe[6][11]),

    .cast_data_o_6_11                               (cast_data_nw_2_pe[6][11]),
    .cast_valid_o_6_11                              (cast_valid_nw_2_pe[6][11]),
    .cast_ready_i_6_11                              (cast_ready_pe_2_nw[6][11]),
    .merge_data_o_6_11                              (merge_data_nw_2_pe[6][11]),
    .merge_valid_o_6_11                             (merge_valid_nw_2_pe[6][11]),
    .merge_ready_i_6_11                             (merge_ready_pe_2_nw[6][11]),
    .gather_data_o_6_11                             (gather_data_nw_2_pe[6][11]),
    .gather_valid_o_6_11                            (gather_valid_nw_2_pe[6][11]),
    .gather_ready_i_6_11                            (gather_ready_pe_2_nw[6][11]),
    .cast_data_i_6_12                               (cast_data_pe_2_nw[6][12]),
    .cast_valid_i_6_12                              (cast_valid_pe_2_nw[6][12]),
    .cast_ready_o_6_12                              (cast_ready_nw_2_pe[6][12]),
    .merge_data_i_6_12                              (merge_data_pe_2_nw[6][12]),
    .merge_valid_i_6_12                             (merge_valid_pe_2_nw[6][12]),
    .merge_ready_o_6_12                             (merge_ready_nw_2_pe[6][12]),
    .gather_data_i_6_12                             (gather_data_pe_2_nw[6][12]),
    .gather_valid_i_6_12                            (gather_valid_pe_2_nw[6][12]),
    .gather_ready_o_6_12                            (gather_ready_nw_2_pe[6][12]),

    .cast_data_o_6_12                               (cast_data_nw_2_pe[6][12]),
    .cast_valid_o_6_12                              (cast_valid_nw_2_pe[6][12]),
    .cast_ready_i_6_12                              (cast_ready_pe_2_nw[6][12]),
    .merge_data_o_6_12                              (merge_data_nw_2_pe[6][12]),
    .merge_valid_o_6_12                             (merge_valid_nw_2_pe[6][12]),
    .merge_ready_i_6_12                             (merge_ready_pe_2_nw[6][12]),
    .gather_data_o_6_12                             (gather_data_nw_2_pe[6][12]),
    .gather_valid_o_6_12                            (gather_valid_nw_2_pe[6][12]),
    .gather_ready_i_6_12                            (gather_ready_pe_2_nw[6][12]),
    .cast_data_i_6_13                               (cast_data_pe_2_nw[6][13]),
    .cast_valid_i_6_13                              (cast_valid_pe_2_nw[6][13]),
    .cast_ready_o_6_13                              (cast_ready_nw_2_pe[6][13]),
    .merge_data_i_6_13                              (merge_data_pe_2_nw[6][13]),
    .merge_valid_i_6_13                             (merge_valid_pe_2_nw[6][13]),
    .merge_ready_o_6_13                             (merge_ready_nw_2_pe[6][13]),
    .gather_data_i_6_13                             (gather_data_pe_2_nw[6][13]),
    .gather_valid_i_6_13                            (gather_valid_pe_2_nw[6][13]),
    .gather_ready_o_6_13                            (gather_ready_nw_2_pe[6][13]),

    .cast_data_o_6_13                               (cast_data_nw_2_pe[6][13]),
    .cast_valid_o_6_13                              (cast_valid_nw_2_pe[6][13]),
    .cast_ready_i_6_13                              (cast_ready_pe_2_nw[6][13]),
    .merge_data_o_6_13                              (merge_data_nw_2_pe[6][13]),
    .merge_valid_o_6_13                             (merge_valid_nw_2_pe[6][13]),
    .merge_ready_i_6_13                             (merge_ready_pe_2_nw[6][13]),
    .gather_data_o_6_13                             (gather_data_nw_2_pe[6][13]),
    .gather_valid_o_6_13                            (gather_valid_nw_2_pe[6][13]),
    .gather_ready_i_6_13                            (gather_ready_pe_2_nw[6][13]),
    .cast_data_i_6_14                               (cast_data_pe_2_nw[6][14]),
    .cast_valid_i_6_14                              (cast_valid_pe_2_nw[6][14]),
    .cast_ready_o_6_14                              (cast_ready_nw_2_pe[6][14]),
    .merge_data_i_6_14                              (merge_data_pe_2_nw[6][14]),
    .merge_valid_i_6_14                             (merge_valid_pe_2_nw[6][14]),
    .merge_ready_o_6_14                             (merge_ready_nw_2_pe[6][14]),
    .gather_data_i_6_14                             (gather_data_pe_2_nw[6][14]),
    .gather_valid_i_6_14                            (gather_valid_pe_2_nw[6][14]),
    .gather_ready_o_6_14                            (gather_ready_nw_2_pe[6][14]),

    .cast_data_o_6_14                               (cast_data_nw_2_pe[6][14]),
    .cast_valid_o_6_14                              (cast_valid_nw_2_pe[6][14]),
    .cast_ready_i_6_14                              (cast_ready_pe_2_nw[6][14]),
    .merge_data_o_6_14                              (merge_data_nw_2_pe[6][14]),
    .merge_valid_o_6_14                             (merge_valid_nw_2_pe[6][14]),
    .merge_ready_i_6_14                             (merge_ready_pe_2_nw[6][14]),
    .gather_data_o_6_14                             (gather_data_nw_2_pe[6][14]),
    .gather_valid_o_6_14                            (gather_valid_nw_2_pe[6][14]),
    .gather_ready_i_6_14                            (gather_ready_pe_2_nw[6][14]),
    .cast_data_i_6_15                               (cast_data_pe_2_nw[6][15]),
    .cast_valid_i_6_15                              (cast_valid_pe_2_nw[6][15]),
    .cast_ready_o_6_15                              (cast_ready_nw_2_pe[6][15]),
    .merge_data_i_6_15                              (merge_data_pe_2_nw[6][15]),
    .merge_valid_i_6_15                             (merge_valid_pe_2_nw[6][15]),
    .merge_ready_o_6_15                             (merge_ready_nw_2_pe[6][15]),
    .gather_data_i_6_15                             (gather_data_pe_2_nw[6][15]),
    .gather_valid_i_6_15                            (gather_valid_pe_2_nw[6][15]),
    .gather_ready_o_6_15                            (gather_ready_nw_2_pe[6][15]),

    .cast_data_o_6_15                               (cast_data_nw_2_pe[6][15]),
    .cast_valid_o_6_15                              (cast_valid_nw_2_pe[6][15]),
    .cast_ready_i_6_15                              (cast_ready_pe_2_nw[6][15]),
    .merge_data_o_6_15                              (merge_data_nw_2_pe[6][15]),
    .merge_valid_o_6_15                             (merge_valid_nw_2_pe[6][15]),
    .merge_ready_i_6_15                             (merge_ready_pe_2_nw[6][15]),
    .gather_data_o_6_15                             (gather_data_nw_2_pe[6][15]),
    .gather_valid_o_6_15                            (gather_valid_nw_2_pe[6][15]),
    .gather_ready_i_6_15                            (gather_ready_pe_2_nw[6][15]),
    .cast_data_i_6_16                               (cast_data_pe_2_nw[6][16]),
    .cast_valid_i_6_16                              (cast_valid_pe_2_nw[6][16]),
    .cast_ready_o_6_16                              (cast_ready_nw_2_pe[6][16]),
    .merge_data_i_6_16                              (merge_data_pe_2_nw[6][16]),
    .merge_valid_i_6_16                             (merge_valid_pe_2_nw[6][16]),
    .merge_ready_o_6_16                             (merge_ready_nw_2_pe[6][16]),
    .gather_data_i_6_16                             (gather_data_pe_2_nw[6][16]),
    .gather_valid_i_6_16                            (gather_valid_pe_2_nw[6][16]),
    .gather_ready_o_6_16                            (gather_ready_nw_2_pe[6][16]),

    .cast_data_o_6_16                               (cast_data_nw_2_pe[6][16]),
    .cast_valid_o_6_16                              (cast_valid_nw_2_pe[6][16]),
    .cast_ready_i_6_16                              (cast_ready_pe_2_nw[6][16]),
    .merge_data_o_6_16                              (merge_data_nw_2_pe[6][16]),
    .merge_valid_o_6_16                             (merge_valid_nw_2_pe[6][16]),
    .merge_ready_i_6_16                             (merge_ready_pe_2_nw[6][16]),
    .gather_data_o_6_16                             (gather_data_nw_2_pe[6][16]),
    .gather_valid_o_6_16                            (gather_valid_nw_2_pe[6][16]),
    .gather_ready_i_6_16                            (gather_ready_pe_2_nw[6][16]),
    .cast_data_i_6_17                               (cast_data_pe_2_nw[6][17]),
    .cast_valid_i_6_17                              (cast_valid_pe_2_nw[6][17]),
    .cast_ready_o_6_17                              (cast_ready_nw_2_pe[6][17]),
    .merge_data_i_6_17                              (merge_data_pe_2_nw[6][17]),
    .merge_valid_i_6_17                             (merge_valid_pe_2_nw[6][17]),
    .merge_ready_o_6_17                             (merge_ready_nw_2_pe[6][17]),
    .gather_data_i_6_17                             (gather_data_pe_2_nw[6][17]),
    .gather_valid_i_6_17                            (gather_valid_pe_2_nw[6][17]),
    .gather_ready_o_6_17                            (gather_ready_nw_2_pe[6][17]),

    .cast_data_o_6_17                               (cast_data_nw_2_pe[6][17]),
    .cast_valid_o_6_17                              (cast_valid_nw_2_pe[6][17]),
    .cast_ready_i_6_17                              (cast_ready_pe_2_nw[6][17]),
    .merge_data_o_6_17                              (merge_data_nw_2_pe[6][17]),
    .merge_valid_o_6_17                             (merge_valid_nw_2_pe[6][17]),
    .merge_ready_i_6_17                             (merge_ready_pe_2_nw[6][17]),
    .gather_data_o_6_17                             (gather_data_nw_2_pe[6][17]),
    .gather_valid_o_6_17                            (gather_valid_nw_2_pe[6][17]),
    .gather_ready_i_6_17                            (gather_ready_pe_2_nw[6][17]),
    .cast_data_i_6_18                               (cast_data_pe_2_nw[6][18]),
    .cast_valid_i_6_18                              (cast_valid_pe_2_nw[6][18]),
    .cast_ready_o_6_18                              (cast_ready_nw_2_pe[6][18]),
    .merge_data_i_6_18                              (merge_data_pe_2_nw[6][18]),
    .merge_valid_i_6_18                             (merge_valid_pe_2_nw[6][18]),
    .merge_ready_o_6_18                             (merge_ready_nw_2_pe[6][18]),
    .gather_data_i_6_18                             (gather_data_pe_2_nw[6][18]),
    .gather_valid_i_6_18                            (gather_valid_pe_2_nw[6][18]),
    .gather_ready_o_6_18                            (gather_ready_nw_2_pe[6][18]),

    .cast_data_o_6_18                               (cast_data_nw_2_pe[6][18]),
    .cast_valid_o_6_18                              (cast_valid_nw_2_pe[6][18]),
    .cast_ready_i_6_18                              (cast_ready_pe_2_nw[6][18]),
    .merge_data_o_6_18                              (merge_data_nw_2_pe[6][18]),
    .merge_valid_o_6_18                             (merge_valid_nw_2_pe[6][18]),
    .merge_ready_i_6_18                             (merge_ready_pe_2_nw[6][18]),
    .gather_data_o_6_18                             (gather_data_nw_2_pe[6][18]),
    .gather_valid_o_6_18                            (gather_valid_nw_2_pe[6][18]),
    .gather_ready_i_6_18                            (gather_ready_pe_2_nw[6][18]),
    .cast_data_i_6_19                               (cast_data_pe_2_nw[6][19]),
    .cast_valid_i_6_19                              (cast_valid_pe_2_nw[6][19]),
    .cast_ready_o_6_19                              (cast_ready_nw_2_pe[6][19]),
    .merge_data_i_6_19                              (merge_data_pe_2_nw[6][19]),
    .merge_valid_i_6_19                             (merge_valid_pe_2_nw[6][19]),
    .merge_ready_o_6_19                             (merge_ready_nw_2_pe[6][19]),
    .gather_data_i_6_19                             (gather_data_pe_2_nw[6][19]),
    .gather_valid_i_6_19                            (gather_valid_pe_2_nw[6][19]),
    .gather_ready_o_6_19                            (gather_ready_nw_2_pe[6][19]),

    .cast_data_o_6_19                               (cast_data_nw_2_pe[6][19]),
    .cast_valid_o_6_19                              (cast_valid_nw_2_pe[6][19]),
    .cast_ready_i_6_19                              (cast_ready_pe_2_nw[6][19]),
    .merge_data_o_6_19                              (merge_data_nw_2_pe[6][19]),
    .merge_valid_o_6_19                             (merge_valid_nw_2_pe[6][19]),
    .merge_ready_i_6_19                             (merge_ready_pe_2_nw[6][19]),
    .gather_data_o_6_19                             (gather_data_nw_2_pe[6][19]),
    .gather_valid_o_6_19                            (gather_valid_nw_2_pe[6][19]),
    .gather_ready_i_6_19                            (gather_ready_pe_2_nw[6][19]),
    .cast_data_i_6_20                               (cast_data_pe_2_nw[6][20]),
    .cast_valid_i_6_20                              (cast_valid_pe_2_nw[6][20]),
    .cast_ready_o_6_20                              (cast_ready_nw_2_pe[6][20]),
    .merge_data_i_6_20                              (merge_data_pe_2_nw[6][20]),
    .merge_valid_i_6_20                             (merge_valid_pe_2_nw[6][20]),
    .merge_ready_o_6_20                             (merge_ready_nw_2_pe[6][20]),
    .gather_data_i_6_20                             (gather_data_pe_2_nw[6][20]),
    .gather_valid_i_6_20                            (gather_valid_pe_2_nw[6][20]),
    .gather_ready_o_6_20                            (gather_ready_nw_2_pe[6][20]),

    .cast_data_o_6_20                               (cast_data_nw_2_pe[6][20]),
    .cast_valid_o_6_20                              (cast_valid_nw_2_pe[6][20]),
    .cast_ready_i_6_20                              (cast_ready_pe_2_nw[6][20]),
    .merge_data_o_6_20                              (merge_data_nw_2_pe[6][20]),
    .merge_valid_o_6_20                             (merge_valid_nw_2_pe[6][20]),
    .merge_ready_i_6_20                             (merge_ready_pe_2_nw[6][20]),
    .gather_data_o_6_20                             (gather_data_nw_2_pe[6][20]),
    .gather_valid_o_6_20                            (gather_valid_nw_2_pe[6][20]),
    .gather_ready_i_6_20                            (gather_ready_pe_2_nw[6][20]),
    .cast_data_i_6_21                               (cast_data_pe_2_nw[6][21]),
    .cast_valid_i_6_21                              (cast_valid_pe_2_nw[6][21]),
    .cast_ready_o_6_21                              (cast_ready_nw_2_pe[6][21]),
    .merge_data_i_6_21                              (merge_data_pe_2_nw[6][21]),
    .merge_valid_i_6_21                             (merge_valid_pe_2_nw[6][21]),
    .merge_ready_o_6_21                             (merge_ready_nw_2_pe[6][21]),
    .gather_data_i_6_21                             (gather_data_pe_2_nw[6][21]),
    .gather_valid_i_6_21                            (gather_valid_pe_2_nw[6][21]),
    .gather_ready_o_6_21                            (gather_ready_nw_2_pe[6][21]),

    .cast_data_o_6_21                               (cast_data_nw_2_pe[6][21]),
    .cast_valid_o_6_21                              (cast_valid_nw_2_pe[6][21]),
    .cast_ready_i_6_21                              (cast_ready_pe_2_nw[6][21]),
    .merge_data_o_6_21                              (merge_data_nw_2_pe[6][21]),
    .merge_valid_o_6_21                             (merge_valid_nw_2_pe[6][21]),
    .merge_ready_i_6_21                             (merge_ready_pe_2_nw[6][21]),
    .gather_data_o_6_21                             (gather_data_nw_2_pe[6][21]),
    .gather_valid_o_6_21                            (gather_valid_nw_2_pe[6][21]),
    .gather_ready_i_6_21                            (gather_ready_pe_2_nw[6][21]),
    .cast_data_i_6_22                               (cast_data_pe_2_nw[6][22]),
    .cast_valid_i_6_22                              (cast_valid_pe_2_nw[6][22]),
    .cast_ready_o_6_22                              (cast_ready_nw_2_pe[6][22]),
    .merge_data_i_6_22                              (merge_data_pe_2_nw[6][22]),
    .merge_valid_i_6_22                             (merge_valid_pe_2_nw[6][22]),
    .merge_ready_o_6_22                             (merge_ready_nw_2_pe[6][22]),
    .gather_data_i_6_22                             (gather_data_pe_2_nw[6][22]),
    .gather_valid_i_6_22                            (gather_valid_pe_2_nw[6][22]),
    .gather_ready_o_6_22                            (gather_ready_nw_2_pe[6][22]),

    .cast_data_o_6_22                               (cast_data_nw_2_pe[6][22]),
    .cast_valid_o_6_22                              (cast_valid_nw_2_pe[6][22]),
    .cast_ready_i_6_22                              (cast_ready_pe_2_nw[6][22]),
    .merge_data_o_6_22                              (merge_data_nw_2_pe[6][22]),
    .merge_valid_o_6_22                             (merge_valid_nw_2_pe[6][22]),
    .merge_ready_i_6_22                             (merge_ready_pe_2_nw[6][22]),
    .gather_data_o_6_22                             (gather_data_nw_2_pe[6][22]),
    .gather_valid_o_6_22                            (gather_valid_nw_2_pe[6][22]),
    .gather_ready_i_6_22                            (gather_ready_pe_2_nw[6][22]),
    .cast_data_i_6_23                               (cast_data_pe_2_nw[6][23]),
    .cast_valid_i_6_23                              (cast_valid_pe_2_nw[6][23]),
    .cast_ready_o_6_23                              (cast_ready_nw_2_pe[6][23]),
    .merge_data_i_6_23                              (merge_data_pe_2_nw[6][23]),
    .merge_valid_i_6_23                             (merge_valid_pe_2_nw[6][23]),
    .merge_ready_o_6_23                             (merge_ready_nw_2_pe[6][23]),
    .gather_data_i_6_23                             (gather_data_pe_2_nw[6][23]),
    .gather_valid_i_6_23                            (gather_valid_pe_2_nw[6][23]),
    .gather_ready_o_6_23                            (gather_ready_nw_2_pe[6][23]),

    .cast_data_o_6_23                               (cast_data_nw_2_pe[6][23]),
    .cast_valid_o_6_23                              (cast_valid_nw_2_pe[6][23]),
    .cast_ready_i_6_23                              (cast_ready_pe_2_nw[6][23]),
    .merge_data_o_6_23                              (merge_data_nw_2_pe[6][23]),
    .merge_valid_o_6_23                             (merge_valid_nw_2_pe[6][23]),
    .merge_ready_i_6_23                             (merge_ready_pe_2_nw[6][23]),
    .gather_data_o_6_23                             (gather_data_nw_2_pe[6][23]),
    .gather_valid_o_6_23                            (gather_valid_nw_2_pe[6][23]),
    .gather_ready_i_6_23                            (gather_ready_pe_2_nw[6][23]),
    .cast_data_i_6_24                               (cast_data_pe_2_nw[6][24]),
    .cast_valid_i_6_24                              (cast_valid_pe_2_nw[6][24]),
    .cast_ready_o_6_24                              (cast_ready_nw_2_pe[6][24]),
    .merge_data_i_6_24                              (merge_data_pe_2_nw[6][24]),
    .merge_valid_i_6_24                             (merge_valid_pe_2_nw[6][24]),
    .merge_ready_o_6_24                             (merge_ready_nw_2_pe[6][24]),
    .gather_data_i_6_24                             (gather_data_pe_2_nw[6][24]),
    .gather_valid_i_6_24                            (gather_valid_pe_2_nw[6][24]),
    .gather_ready_o_6_24                            (gather_ready_nw_2_pe[6][24]),

    .cast_data_o_6_24                               (cast_data_nw_2_pe[6][24]),
    .cast_valid_o_6_24                              (cast_valid_nw_2_pe[6][24]),
    .cast_ready_i_6_24                              (cast_ready_pe_2_nw[6][24]),
    .merge_data_o_6_24                              (merge_data_nw_2_pe[6][24]),
    .merge_valid_o_6_24                             (merge_valid_nw_2_pe[6][24]),
    .merge_ready_i_6_24                             (merge_ready_pe_2_nw[6][24]),
    .gather_data_o_6_24                             (gather_data_nw_2_pe[6][24]),
    .gather_valid_o_6_24                            (gather_valid_nw_2_pe[6][24]),
    .gather_ready_i_6_24                            (gather_ready_pe_2_nw[6][24]),
    .cast_data_i_7_0                               (cast_data_pe_2_nw[7][0]),
    .cast_valid_i_7_0                              (cast_valid_pe_2_nw[7][0]),
    .cast_ready_o_7_0                              (cast_ready_nw_2_pe[7][0]),
    .merge_data_i_7_0                              (merge_data_pe_2_nw[7][0]),
    .merge_valid_i_7_0                             (merge_valid_pe_2_nw[7][0]),
    .merge_ready_o_7_0                             (merge_ready_nw_2_pe[7][0]),
    .gather_data_i_7_0                             (gather_data_pe_2_nw[7][0]),
    .gather_valid_i_7_0                            (gather_valid_pe_2_nw[7][0]),
    .gather_ready_o_7_0                            (gather_ready_nw_2_pe[7][0]),

    .cast_data_o_7_0                               (cast_data_nw_2_pe[7][0]),
    .cast_valid_o_7_0                              (cast_valid_nw_2_pe[7][0]),
    .cast_ready_i_7_0                              (cast_ready_pe_2_nw[7][0]),
    .merge_data_o_7_0                              (merge_data_nw_2_pe[7][0]),
    .merge_valid_o_7_0                             (merge_valid_nw_2_pe[7][0]),
    .merge_ready_i_7_0                             (merge_ready_pe_2_nw[7][0]),
    .gather_data_o_7_0                             (gather_data_nw_2_pe[7][0]),
    .gather_valid_o_7_0                            (gather_valid_nw_2_pe[7][0]),
    .gather_ready_i_7_0                            (gather_ready_pe_2_nw[7][0]),
    .cast_data_i_7_1                               (cast_data_pe_2_nw[7][1]),
    .cast_valid_i_7_1                              (cast_valid_pe_2_nw[7][1]),
    .cast_ready_o_7_1                              (cast_ready_nw_2_pe[7][1]),
    .merge_data_i_7_1                              (merge_data_pe_2_nw[7][1]),
    .merge_valid_i_7_1                             (merge_valid_pe_2_nw[7][1]),
    .merge_ready_o_7_1                             (merge_ready_nw_2_pe[7][1]),
    .gather_data_i_7_1                             (gather_data_pe_2_nw[7][1]),
    .gather_valid_i_7_1                            (gather_valid_pe_2_nw[7][1]),
    .gather_ready_o_7_1                            (gather_ready_nw_2_pe[7][1]),

    .cast_data_o_7_1                               (cast_data_nw_2_pe[7][1]),
    .cast_valid_o_7_1                              (cast_valid_nw_2_pe[7][1]),
    .cast_ready_i_7_1                              (cast_ready_pe_2_nw[7][1]),
    .merge_data_o_7_1                              (merge_data_nw_2_pe[7][1]),
    .merge_valid_o_7_1                             (merge_valid_nw_2_pe[7][1]),
    .merge_ready_i_7_1                             (merge_ready_pe_2_nw[7][1]),
    .gather_data_o_7_1                             (gather_data_nw_2_pe[7][1]),
    .gather_valid_o_7_1                            (gather_valid_nw_2_pe[7][1]),
    .gather_ready_i_7_1                            (gather_ready_pe_2_nw[7][1]),
    .cast_data_i_7_2                               (cast_data_pe_2_nw[7][2]),
    .cast_valid_i_7_2                              (cast_valid_pe_2_nw[7][2]),
    .cast_ready_o_7_2                              (cast_ready_nw_2_pe[7][2]),
    .merge_data_i_7_2                              (merge_data_pe_2_nw[7][2]),
    .merge_valid_i_7_2                             (merge_valid_pe_2_nw[7][2]),
    .merge_ready_o_7_2                             (merge_ready_nw_2_pe[7][2]),
    .gather_data_i_7_2                             (gather_data_pe_2_nw[7][2]),
    .gather_valid_i_7_2                            (gather_valid_pe_2_nw[7][2]),
    .gather_ready_o_7_2                            (gather_ready_nw_2_pe[7][2]),

    .cast_data_o_7_2                               (cast_data_nw_2_pe[7][2]),
    .cast_valid_o_7_2                              (cast_valid_nw_2_pe[7][2]),
    .cast_ready_i_7_2                              (cast_ready_pe_2_nw[7][2]),
    .merge_data_o_7_2                              (merge_data_nw_2_pe[7][2]),
    .merge_valid_o_7_2                             (merge_valid_nw_2_pe[7][2]),
    .merge_ready_i_7_2                             (merge_ready_pe_2_nw[7][2]),
    .gather_data_o_7_2                             (gather_data_nw_2_pe[7][2]),
    .gather_valid_o_7_2                            (gather_valid_nw_2_pe[7][2]),
    .gather_ready_i_7_2                            (gather_ready_pe_2_nw[7][2]),
    .cast_data_i_7_3                               (cast_data_pe_2_nw[7][3]),
    .cast_valid_i_7_3                              (cast_valid_pe_2_nw[7][3]),
    .cast_ready_o_7_3                              (cast_ready_nw_2_pe[7][3]),
    .merge_data_i_7_3                              (merge_data_pe_2_nw[7][3]),
    .merge_valid_i_7_3                             (merge_valid_pe_2_nw[7][3]),
    .merge_ready_o_7_3                             (merge_ready_nw_2_pe[7][3]),
    .gather_data_i_7_3                             (gather_data_pe_2_nw[7][3]),
    .gather_valid_i_7_3                            (gather_valid_pe_2_nw[7][3]),
    .gather_ready_o_7_3                            (gather_ready_nw_2_pe[7][3]),

    .cast_data_o_7_3                               (cast_data_nw_2_pe[7][3]),
    .cast_valid_o_7_3                              (cast_valid_nw_2_pe[7][3]),
    .cast_ready_i_7_3                              (cast_ready_pe_2_nw[7][3]),
    .merge_data_o_7_3                              (merge_data_nw_2_pe[7][3]),
    .merge_valid_o_7_3                             (merge_valid_nw_2_pe[7][3]),
    .merge_ready_i_7_3                             (merge_ready_pe_2_nw[7][3]),
    .gather_data_o_7_3                             (gather_data_nw_2_pe[7][3]),
    .gather_valid_o_7_3                            (gather_valid_nw_2_pe[7][3]),
    .gather_ready_i_7_3                            (gather_ready_pe_2_nw[7][3]),
    .cast_data_i_7_4                               (cast_data_pe_2_nw[7][4]),
    .cast_valid_i_7_4                              (cast_valid_pe_2_nw[7][4]),
    .cast_ready_o_7_4                              (cast_ready_nw_2_pe[7][4]),
    .merge_data_i_7_4                              (merge_data_pe_2_nw[7][4]),
    .merge_valid_i_7_4                             (merge_valid_pe_2_nw[7][4]),
    .merge_ready_o_7_4                             (merge_ready_nw_2_pe[7][4]),
    .gather_data_i_7_4                             (gather_data_pe_2_nw[7][4]),
    .gather_valid_i_7_4                            (gather_valid_pe_2_nw[7][4]),
    .gather_ready_o_7_4                            (gather_ready_nw_2_pe[7][4]),

    .cast_data_o_7_4                               (cast_data_nw_2_pe[7][4]),
    .cast_valid_o_7_4                              (cast_valid_nw_2_pe[7][4]),
    .cast_ready_i_7_4                              (cast_ready_pe_2_nw[7][4]),
    .merge_data_o_7_4                              (merge_data_nw_2_pe[7][4]),
    .merge_valid_o_7_4                             (merge_valid_nw_2_pe[7][4]),
    .merge_ready_i_7_4                             (merge_ready_pe_2_nw[7][4]),
    .gather_data_o_7_4                             (gather_data_nw_2_pe[7][4]),
    .gather_valid_o_7_4                            (gather_valid_nw_2_pe[7][4]),
    .gather_ready_i_7_4                            (gather_ready_pe_2_nw[7][4]),
    .cast_data_i_7_5                               (cast_data_pe_2_nw[7][5]),
    .cast_valid_i_7_5                              (cast_valid_pe_2_nw[7][5]),
    .cast_ready_o_7_5                              (cast_ready_nw_2_pe[7][5]),
    .merge_data_i_7_5                              (merge_data_pe_2_nw[7][5]),
    .merge_valid_i_7_5                             (merge_valid_pe_2_nw[7][5]),
    .merge_ready_o_7_5                             (merge_ready_nw_2_pe[7][5]),
    .gather_data_i_7_5                             (gather_data_pe_2_nw[7][5]),
    .gather_valid_i_7_5                            (gather_valid_pe_2_nw[7][5]),
    .gather_ready_o_7_5                            (gather_ready_nw_2_pe[7][5]),

    .cast_data_o_7_5                               (cast_data_nw_2_pe[7][5]),
    .cast_valid_o_7_5                              (cast_valid_nw_2_pe[7][5]),
    .cast_ready_i_7_5                              (cast_ready_pe_2_nw[7][5]),
    .merge_data_o_7_5                              (merge_data_nw_2_pe[7][5]),
    .merge_valid_o_7_5                             (merge_valid_nw_2_pe[7][5]),
    .merge_ready_i_7_5                             (merge_ready_pe_2_nw[7][5]),
    .gather_data_o_7_5                             (gather_data_nw_2_pe[7][5]),
    .gather_valid_o_7_5                            (gather_valid_nw_2_pe[7][5]),
    .gather_ready_i_7_5                            (gather_ready_pe_2_nw[7][5]),
    .cast_data_i_7_6                               (cast_data_pe_2_nw[7][6]),
    .cast_valid_i_7_6                              (cast_valid_pe_2_nw[7][6]),
    .cast_ready_o_7_6                              (cast_ready_nw_2_pe[7][6]),
    .merge_data_i_7_6                              (merge_data_pe_2_nw[7][6]),
    .merge_valid_i_7_6                             (merge_valid_pe_2_nw[7][6]),
    .merge_ready_o_7_6                             (merge_ready_nw_2_pe[7][6]),
    .gather_data_i_7_6                             (gather_data_pe_2_nw[7][6]),
    .gather_valid_i_7_6                            (gather_valid_pe_2_nw[7][6]),
    .gather_ready_o_7_6                            (gather_ready_nw_2_pe[7][6]),

    .cast_data_o_7_6                               (cast_data_nw_2_pe[7][6]),
    .cast_valid_o_7_6                              (cast_valid_nw_2_pe[7][6]),
    .cast_ready_i_7_6                              (cast_ready_pe_2_nw[7][6]),
    .merge_data_o_7_6                              (merge_data_nw_2_pe[7][6]),
    .merge_valid_o_7_6                             (merge_valid_nw_2_pe[7][6]),
    .merge_ready_i_7_6                             (merge_ready_pe_2_nw[7][6]),
    .gather_data_o_7_6                             (gather_data_nw_2_pe[7][6]),
    .gather_valid_o_7_6                            (gather_valid_nw_2_pe[7][6]),
    .gather_ready_i_7_6                            (gather_ready_pe_2_nw[7][6]),
    .cast_data_i_7_7                               (cast_data_pe_2_nw[7][7]),
    .cast_valid_i_7_7                              (cast_valid_pe_2_nw[7][7]),
    .cast_ready_o_7_7                              (cast_ready_nw_2_pe[7][7]),
    .merge_data_i_7_7                              (merge_data_pe_2_nw[7][7]),
    .merge_valid_i_7_7                             (merge_valid_pe_2_nw[7][7]),
    .merge_ready_o_7_7                             (merge_ready_nw_2_pe[7][7]),
    .gather_data_i_7_7                             (gather_data_pe_2_nw[7][7]),
    .gather_valid_i_7_7                            (gather_valid_pe_2_nw[7][7]),
    .gather_ready_o_7_7                            (gather_ready_nw_2_pe[7][7]),

    .cast_data_o_7_7                               (cast_data_nw_2_pe[7][7]),
    .cast_valid_o_7_7                              (cast_valid_nw_2_pe[7][7]),
    .cast_ready_i_7_7                              (cast_ready_pe_2_nw[7][7]),
    .merge_data_o_7_7                              (merge_data_nw_2_pe[7][7]),
    .merge_valid_o_7_7                             (merge_valid_nw_2_pe[7][7]),
    .merge_ready_i_7_7                             (merge_ready_pe_2_nw[7][7]),
    .gather_data_o_7_7                             (gather_data_nw_2_pe[7][7]),
    .gather_valid_o_7_7                            (gather_valid_nw_2_pe[7][7]),
    .gather_ready_i_7_7                            (gather_ready_pe_2_nw[7][7]),
    .cast_data_i_7_8                               (cast_data_pe_2_nw[7][8]),
    .cast_valid_i_7_8                              (cast_valid_pe_2_nw[7][8]),
    .cast_ready_o_7_8                              (cast_ready_nw_2_pe[7][8]),
    .merge_data_i_7_8                              (merge_data_pe_2_nw[7][8]),
    .merge_valid_i_7_8                             (merge_valid_pe_2_nw[7][8]),
    .merge_ready_o_7_8                             (merge_ready_nw_2_pe[7][8]),
    .gather_data_i_7_8                             (gather_data_pe_2_nw[7][8]),
    .gather_valid_i_7_8                            (gather_valid_pe_2_nw[7][8]),
    .gather_ready_o_7_8                            (gather_ready_nw_2_pe[7][8]),

    .cast_data_o_7_8                               (cast_data_nw_2_pe[7][8]),
    .cast_valid_o_7_8                              (cast_valid_nw_2_pe[7][8]),
    .cast_ready_i_7_8                              (cast_ready_pe_2_nw[7][8]),
    .merge_data_o_7_8                              (merge_data_nw_2_pe[7][8]),
    .merge_valid_o_7_8                             (merge_valid_nw_2_pe[7][8]),
    .merge_ready_i_7_8                             (merge_ready_pe_2_nw[7][8]),
    .gather_data_o_7_8                             (gather_data_nw_2_pe[7][8]),
    .gather_valid_o_7_8                            (gather_valid_nw_2_pe[7][8]),
    .gather_ready_i_7_8                            (gather_ready_pe_2_nw[7][8]),
    .cast_data_i_7_9                               (cast_data_pe_2_nw[7][9]),
    .cast_valid_i_7_9                              (cast_valid_pe_2_nw[7][9]),
    .cast_ready_o_7_9                              (cast_ready_nw_2_pe[7][9]),
    .merge_data_i_7_9                              (merge_data_pe_2_nw[7][9]),
    .merge_valid_i_7_9                             (merge_valid_pe_2_nw[7][9]),
    .merge_ready_o_7_9                             (merge_ready_nw_2_pe[7][9]),
    .gather_data_i_7_9                             (gather_data_pe_2_nw[7][9]),
    .gather_valid_i_7_9                            (gather_valid_pe_2_nw[7][9]),
    .gather_ready_o_7_9                            (gather_ready_nw_2_pe[7][9]),

    .cast_data_o_7_9                               (cast_data_nw_2_pe[7][9]),
    .cast_valid_o_7_9                              (cast_valid_nw_2_pe[7][9]),
    .cast_ready_i_7_9                              (cast_ready_pe_2_nw[7][9]),
    .merge_data_o_7_9                              (merge_data_nw_2_pe[7][9]),
    .merge_valid_o_7_9                             (merge_valid_nw_2_pe[7][9]),
    .merge_ready_i_7_9                             (merge_ready_pe_2_nw[7][9]),
    .gather_data_o_7_9                             (gather_data_nw_2_pe[7][9]),
    .gather_valid_o_7_9                            (gather_valid_nw_2_pe[7][9]),
    .gather_ready_i_7_9                            (gather_ready_pe_2_nw[7][9]),
    .cast_data_i_7_10                               (cast_data_pe_2_nw[7][10]),
    .cast_valid_i_7_10                              (cast_valid_pe_2_nw[7][10]),
    .cast_ready_o_7_10                              (cast_ready_nw_2_pe[7][10]),
    .merge_data_i_7_10                              (merge_data_pe_2_nw[7][10]),
    .merge_valid_i_7_10                             (merge_valid_pe_2_nw[7][10]),
    .merge_ready_o_7_10                             (merge_ready_nw_2_pe[7][10]),
    .gather_data_i_7_10                             (gather_data_pe_2_nw[7][10]),
    .gather_valid_i_7_10                            (gather_valid_pe_2_nw[7][10]),
    .gather_ready_o_7_10                            (gather_ready_nw_2_pe[7][10]),

    .cast_data_o_7_10                               (cast_data_nw_2_pe[7][10]),
    .cast_valid_o_7_10                              (cast_valid_nw_2_pe[7][10]),
    .cast_ready_i_7_10                              (cast_ready_pe_2_nw[7][10]),
    .merge_data_o_7_10                              (merge_data_nw_2_pe[7][10]),
    .merge_valid_o_7_10                             (merge_valid_nw_2_pe[7][10]),
    .merge_ready_i_7_10                             (merge_ready_pe_2_nw[7][10]),
    .gather_data_o_7_10                             (gather_data_nw_2_pe[7][10]),
    .gather_valid_o_7_10                            (gather_valid_nw_2_pe[7][10]),
    .gather_ready_i_7_10                            (gather_ready_pe_2_nw[7][10]),
    .cast_data_i_7_11                               (cast_data_pe_2_nw[7][11]),
    .cast_valid_i_7_11                              (cast_valid_pe_2_nw[7][11]),
    .cast_ready_o_7_11                              (cast_ready_nw_2_pe[7][11]),
    .merge_data_i_7_11                              (merge_data_pe_2_nw[7][11]),
    .merge_valid_i_7_11                             (merge_valid_pe_2_nw[7][11]),
    .merge_ready_o_7_11                             (merge_ready_nw_2_pe[7][11]),
    .gather_data_i_7_11                             (gather_data_pe_2_nw[7][11]),
    .gather_valid_i_7_11                            (gather_valid_pe_2_nw[7][11]),
    .gather_ready_o_7_11                            (gather_ready_nw_2_pe[7][11]),

    .cast_data_o_7_11                               (cast_data_nw_2_pe[7][11]),
    .cast_valid_o_7_11                              (cast_valid_nw_2_pe[7][11]),
    .cast_ready_i_7_11                              (cast_ready_pe_2_nw[7][11]),
    .merge_data_o_7_11                              (merge_data_nw_2_pe[7][11]),
    .merge_valid_o_7_11                             (merge_valid_nw_2_pe[7][11]),
    .merge_ready_i_7_11                             (merge_ready_pe_2_nw[7][11]),
    .gather_data_o_7_11                             (gather_data_nw_2_pe[7][11]),
    .gather_valid_o_7_11                            (gather_valid_nw_2_pe[7][11]),
    .gather_ready_i_7_11                            (gather_ready_pe_2_nw[7][11]),
    .cast_data_i_7_12                               (cast_data_pe_2_nw[7][12]),
    .cast_valid_i_7_12                              (cast_valid_pe_2_nw[7][12]),
    .cast_ready_o_7_12                              (cast_ready_nw_2_pe[7][12]),
    .merge_data_i_7_12                              (merge_data_pe_2_nw[7][12]),
    .merge_valid_i_7_12                             (merge_valid_pe_2_nw[7][12]),
    .merge_ready_o_7_12                             (merge_ready_nw_2_pe[7][12]),
    .gather_data_i_7_12                             (gather_data_pe_2_nw[7][12]),
    .gather_valid_i_7_12                            (gather_valid_pe_2_nw[7][12]),
    .gather_ready_o_7_12                            (gather_ready_nw_2_pe[7][12]),

    .cast_data_o_7_12                               (cast_data_nw_2_pe[7][12]),
    .cast_valid_o_7_12                              (cast_valid_nw_2_pe[7][12]),
    .cast_ready_i_7_12                              (cast_ready_pe_2_nw[7][12]),
    .merge_data_o_7_12                              (merge_data_nw_2_pe[7][12]),
    .merge_valid_o_7_12                             (merge_valid_nw_2_pe[7][12]),
    .merge_ready_i_7_12                             (merge_ready_pe_2_nw[7][12]),
    .gather_data_o_7_12                             (gather_data_nw_2_pe[7][12]),
    .gather_valid_o_7_12                            (gather_valid_nw_2_pe[7][12]),
    .gather_ready_i_7_12                            (gather_ready_pe_2_nw[7][12]),
    .cast_data_i_7_13                               (cast_data_pe_2_nw[7][13]),
    .cast_valid_i_7_13                              (cast_valid_pe_2_nw[7][13]),
    .cast_ready_o_7_13                              (cast_ready_nw_2_pe[7][13]),
    .merge_data_i_7_13                              (merge_data_pe_2_nw[7][13]),
    .merge_valid_i_7_13                             (merge_valid_pe_2_nw[7][13]),
    .merge_ready_o_7_13                             (merge_ready_nw_2_pe[7][13]),
    .gather_data_i_7_13                             (gather_data_pe_2_nw[7][13]),
    .gather_valid_i_7_13                            (gather_valid_pe_2_nw[7][13]),
    .gather_ready_o_7_13                            (gather_ready_nw_2_pe[7][13]),

    .cast_data_o_7_13                               (cast_data_nw_2_pe[7][13]),
    .cast_valid_o_7_13                              (cast_valid_nw_2_pe[7][13]),
    .cast_ready_i_7_13                              (cast_ready_pe_2_nw[7][13]),
    .merge_data_o_7_13                              (merge_data_nw_2_pe[7][13]),
    .merge_valid_o_7_13                             (merge_valid_nw_2_pe[7][13]),
    .merge_ready_i_7_13                             (merge_ready_pe_2_nw[7][13]),
    .gather_data_o_7_13                             (gather_data_nw_2_pe[7][13]),
    .gather_valid_o_7_13                            (gather_valid_nw_2_pe[7][13]),
    .gather_ready_i_7_13                            (gather_ready_pe_2_nw[7][13]),
    .cast_data_i_7_14                               (cast_data_pe_2_nw[7][14]),
    .cast_valid_i_7_14                              (cast_valid_pe_2_nw[7][14]),
    .cast_ready_o_7_14                              (cast_ready_nw_2_pe[7][14]),
    .merge_data_i_7_14                              (merge_data_pe_2_nw[7][14]),
    .merge_valid_i_7_14                             (merge_valid_pe_2_nw[7][14]),
    .merge_ready_o_7_14                             (merge_ready_nw_2_pe[7][14]),
    .gather_data_i_7_14                             (gather_data_pe_2_nw[7][14]),
    .gather_valid_i_7_14                            (gather_valid_pe_2_nw[7][14]),
    .gather_ready_o_7_14                            (gather_ready_nw_2_pe[7][14]),

    .cast_data_o_7_14                               (cast_data_nw_2_pe[7][14]),
    .cast_valid_o_7_14                              (cast_valid_nw_2_pe[7][14]),
    .cast_ready_i_7_14                              (cast_ready_pe_2_nw[7][14]),
    .merge_data_o_7_14                              (merge_data_nw_2_pe[7][14]),
    .merge_valid_o_7_14                             (merge_valid_nw_2_pe[7][14]),
    .merge_ready_i_7_14                             (merge_ready_pe_2_nw[7][14]),
    .gather_data_o_7_14                             (gather_data_nw_2_pe[7][14]),
    .gather_valid_o_7_14                            (gather_valid_nw_2_pe[7][14]),
    .gather_ready_i_7_14                            (gather_ready_pe_2_nw[7][14]),
    .cast_data_i_7_15                               (cast_data_pe_2_nw[7][15]),
    .cast_valid_i_7_15                              (cast_valid_pe_2_nw[7][15]),
    .cast_ready_o_7_15                              (cast_ready_nw_2_pe[7][15]),
    .merge_data_i_7_15                              (merge_data_pe_2_nw[7][15]),
    .merge_valid_i_7_15                             (merge_valid_pe_2_nw[7][15]),
    .merge_ready_o_7_15                             (merge_ready_nw_2_pe[7][15]),
    .gather_data_i_7_15                             (gather_data_pe_2_nw[7][15]),
    .gather_valid_i_7_15                            (gather_valid_pe_2_nw[7][15]),
    .gather_ready_o_7_15                            (gather_ready_nw_2_pe[7][15]),

    .cast_data_o_7_15                               (cast_data_nw_2_pe[7][15]),
    .cast_valid_o_7_15                              (cast_valid_nw_2_pe[7][15]),
    .cast_ready_i_7_15                              (cast_ready_pe_2_nw[7][15]),
    .merge_data_o_7_15                              (merge_data_nw_2_pe[7][15]),
    .merge_valid_o_7_15                             (merge_valid_nw_2_pe[7][15]),
    .merge_ready_i_7_15                             (merge_ready_pe_2_nw[7][15]),
    .gather_data_o_7_15                             (gather_data_nw_2_pe[7][15]),
    .gather_valid_o_7_15                            (gather_valid_nw_2_pe[7][15]),
    .gather_ready_i_7_15                            (gather_ready_pe_2_nw[7][15]),
    .cast_data_i_7_16                               (cast_data_pe_2_nw[7][16]),
    .cast_valid_i_7_16                              (cast_valid_pe_2_nw[7][16]),
    .cast_ready_o_7_16                              (cast_ready_nw_2_pe[7][16]),
    .merge_data_i_7_16                              (merge_data_pe_2_nw[7][16]),
    .merge_valid_i_7_16                             (merge_valid_pe_2_nw[7][16]),
    .merge_ready_o_7_16                             (merge_ready_nw_2_pe[7][16]),
    .gather_data_i_7_16                             (gather_data_pe_2_nw[7][16]),
    .gather_valid_i_7_16                            (gather_valid_pe_2_nw[7][16]),
    .gather_ready_o_7_16                            (gather_ready_nw_2_pe[7][16]),

    .cast_data_o_7_16                               (cast_data_nw_2_pe[7][16]),
    .cast_valid_o_7_16                              (cast_valid_nw_2_pe[7][16]),
    .cast_ready_i_7_16                              (cast_ready_pe_2_nw[7][16]),
    .merge_data_o_7_16                              (merge_data_nw_2_pe[7][16]),
    .merge_valid_o_7_16                             (merge_valid_nw_2_pe[7][16]),
    .merge_ready_i_7_16                             (merge_ready_pe_2_nw[7][16]),
    .gather_data_o_7_16                             (gather_data_nw_2_pe[7][16]),
    .gather_valid_o_7_16                            (gather_valid_nw_2_pe[7][16]),
    .gather_ready_i_7_16                            (gather_ready_pe_2_nw[7][16]),
    .cast_data_i_7_17                               (cast_data_pe_2_nw[7][17]),
    .cast_valid_i_7_17                              (cast_valid_pe_2_nw[7][17]),
    .cast_ready_o_7_17                              (cast_ready_nw_2_pe[7][17]),
    .merge_data_i_7_17                              (merge_data_pe_2_nw[7][17]),
    .merge_valid_i_7_17                             (merge_valid_pe_2_nw[7][17]),
    .merge_ready_o_7_17                             (merge_ready_nw_2_pe[7][17]),
    .gather_data_i_7_17                             (gather_data_pe_2_nw[7][17]),
    .gather_valid_i_7_17                            (gather_valid_pe_2_nw[7][17]),
    .gather_ready_o_7_17                            (gather_ready_nw_2_pe[7][17]),

    .cast_data_o_7_17                               (cast_data_nw_2_pe[7][17]),
    .cast_valid_o_7_17                              (cast_valid_nw_2_pe[7][17]),
    .cast_ready_i_7_17                              (cast_ready_pe_2_nw[7][17]),
    .merge_data_o_7_17                              (merge_data_nw_2_pe[7][17]),
    .merge_valid_o_7_17                             (merge_valid_nw_2_pe[7][17]),
    .merge_ready_i_7_17                             (merge_ready_pe_2_nw[7][17]),
    .gather_data_o_7_17                             (gather_data_nw_2_pe[7][17]),
    .gather_valid_o_7_17                            (gather_valid_nw_2_pe[7][17]),
    .gather_ready_i_7_17                            (gather_ready_pe_2_nw[7][17]),
    .cast_data_i_7_18                               (cast_data_pe_2_nw[7][18]),
    .cast_valid_i_7_18                              (cast_valid_pe_2_nw[7][18]),
    .cast_ready_o_7_18                              (cast_ready_nw_2_pe[7][18]),
    .merge_data_i_7_18                              (merge_data_pe_2_nw[7][18]),
    .merge_valid_i_7_18                             (merge_valid_pe_2_nw[7][18]),
    .merge_ready_o_7_18                             (merge_ready_nw_2_pe[7][18]),
    .gather_data_i_7_18                             (gather_data_pe_2_nw[7][18]),
    .gather_valid_i_7_18                            (gather_valid_pe_2_nw[7][18]),
    .gather_ready_o_7_18                            (gather_ready_nw_2_pe[7][18]),

    .cast_data_o_7_18                               (cast_data_nw_2_pe[7][18]),
    .cast_valid_o_7_18                              (cast_valid_nw_2_pe[7][18]),
    .cast_ready_i_7_18                              (cast_ready_pe_2_nw[7][18]),
    .merge_data_o_7_18                              (merge_data_nw_2_pe[7][18]),
    .merge_valid_o_7_18                             (merge_valid_nw_2_pe[7][18]),
    .merge_ready_i_7_18                             (merge_ready_pe_2_nw[7][18]),
    .gather_data_o_7_18                             (gather_data_nw_2_pe[7][18]),
    .gather_valid_o_7_18                            (gather_valid_nw_2_pe[7][18]),
    .gather_ready_i_7_18                            (gather_ready_pe_2_nw[7][18]),
    .cast_data_i_7_19                               (cast_data_pe_2_nw[7][19]),
    .cast_valid_i_7_19                              (cast_valid_pe_2_nw[7][19]),
    .cast_ready_o_7_19                              (cast_ready_nw_2_pe[7][19]),
    .merge_data_i_7_19                              (merge_data_pe_2_nw[7][19]),
    .merge_valid_i_7_19                             (merge_valid_pe_2_nw[7][19]),
    .merge_ready_o_7_19                             (merge_ready_nw_2_pe[7][19]),
    .gather_data_i_7_19                             (gather_data_pe_2_nw[7][19]),
    .gather_valid_i_7_19                            (gather_valid_pe_2_nw[7][19]),
    .gather_ready_o_7_19                            (gather_ready_nw_2_pe[7][19]),

    .cast_data_o_7_19                               (cast_data_nw_2_pe[7][19]),
    .cast_valid_o_7_19                              (cast_valid_nw_2_pe[7][19]),
    .cast_ready_i_7_19                              (cast_ready_pe_2_nw[7][19]),
    .merge_data_o_7_19                              (merge_data_nw_2_pe[7][19]),
    .merge_valid_o_7_19                             (merge_valid_nw_2_pe[7][19]),
    .merge_ready_i_7_19                             (merge_ready_pe_2_nw[7][19]),
    .gather_data_o_7_19                             (gather_data_nw_2_pe[7][19]),
    .gather_valid_o_7_19                            (gather_valid_nw_2_pe[7][19]),
    .gather_ready_i_7_19                            (gather_ready_pe_2_nw[7][19]),
    .cast_data_i_7_20                               (cast_data_pe_2_nw[7][20]),
    .cast_valid_i_7_20                              (cast_valid_pe_2_nw[7][20]),
    .cast_ready_o_7_20                              (cast_ready_nw_2_pe[7][20]),
    .merge_data_i_7_20                              (merge_data_pe_2_nw[7][20]),
    .merge_valid_i_7_20                             (merge_valid_pe_2_nw[7][20]),
    .merge_ready_o_7_20                             (merge_ready_nw_2_pe[7][20]),
    .gather_data_i_7_20                             (gather_data_pe_2_nw[7][20]),
    .gather_valid_i_7_20                            (gather_valid_pe_2_nw[7][20]),
    .gather_ready_o_7_20                            (gather_ready_nw_2_pe[7][20]),

    .cast_data_o_7_20                               (cast_data_nw_2_pe[7][20]),
    .cast_valid_o_7_20                              (cast_valid_nw_2_pe[7][20]),
    .cast_ready_i_7_20                              (cast_ready_pe_2_nw[7][20]),
    .merge_data_o_7_20                              (merge_data_nw_2_pe[7][20]),
    .merge_valid_o_7_20                             (merge_valid_nw_2_pe[7][20]),
    .merge_ready_i_7_20                             (merge_ready_pe_2_nw[7][20]),
    .gather_data_o_7_20                             (gather_data_nw_2_pe[7][20]),
    .gather_valid_o_7_20                            (gather_valid_nw_2_pe[7][20]),
    .gather_ready_i_7_20                            (gather_ready_pe_2_nw[7][20]),
    .cast_data_i_7_21                               (cast_data_pe_2_nw[7][21]),
    .cast_valid_i_7_21                              (cast_valid_pe_2_nw[7][21]),
    .cast_ready_o_7_21                              (cast_ready_nw_2_pe[7][21]),
    .merge_data_i_7_21                              (merge_data_pe_2_nw[7][21]),
    .merge_valid_i_7_21                             (merge_valid_pe_2_nw[7][21]),
    .merge_ready_o_7_21                             (merge_ready_nw_2_pe[7][21]),
    .gather_data_i_7_21                             (gather_data_pe_2_nw[7][21]),
    .gather_valid_i_7_21                            (gather_valid_pe_2_nw[7][21]),
    .gather_ready_o_7_21                            (gather_ready_nw_2_pe[7][21]),

    .cast_data_o_7_21                               (cast_data_nw_2_pe[7][21]),
    .cast_valid_o_7_21                              (cast_valid_nw_2_pe[7][21]),
    .cast_ready_i_7_21                              (cast_ready_pe_2_nw[7][21]),
    .merge_data_o_7_21                              (merge_data_nw_2_pe[7][21]),
    .merge_valid_o_7_21                             (merge_valid_nw_2_pe[7][21]),
    .merge_ready_i_7_21                             (merge_ready_pe_2_nw[7][21]),
    .gather_data_o_7_21                             (gather_data_nw_2_pe[7][21]),
    .gather_valid_o_7_21                            (gather_valid_nw_2_pe[7][21]),
    .gather_ready_i_7_21                            (gather_ready_pe_2_nw[7][21]),
    .cast_data_i_7_22                               (cast_data_pe_2_nw[7][22]),
    .cast_valid_i_7_22                              (cast_valid_pe_2_nw[7][22]),
    .cast_ready_o_7_22                              (cast_ready_nw_2_pe[7][22]),
    .merge_data_i_7_22                              (merge_data_pe_2_nw[7][22]),
    .merge_valid_i_7_22                             (merge_valid_pe_2_nw[7][22]),
    .merge_ready_o_7_22                             (merge_ready_nw_2_pe[7][22]),
    .gather_data_i_7_22                             (gather_data_pe_2_nw[7][22]),
    .gather_valid_i_7_22                            (gather_valid_pe_2_nw[7][22]),
    .gather_ready_o_7_22                            (gather_ready_nw_2_pe[7][22]),

    .cast_data_o_7_22                               (cast_data_nw_2_pe[7][22]),
    .cast_valid_o_7_22                              (cast_valid_nw_2_pe[7][22]),
    .cast_ready_i_7_22                              (cast_ready_pe_2_nw[7][22]),
    .merge_data_o_7_22                              (merge_data_nw_2_pe[7][22]),
    .merge_valid_o_7_22                             (merge_valid_nw_2_pe[7][22]),
    .merge_ready_i_7_22                             (merge_ready_pe_2_nw[7][22]),
    .gather_data_o_7_22                             (gather_data_nw_2_pe[7][22]),
    .gather_valid_o_7_22                            (gather_valid_nw_2_pe[7][22]),
    .gather_ready_i_7_22                            (gather_ready_pe_2_nw[7][22]),
    .cast_data_i_7_23                               (cast_data_pe_2_nw[7][23]),
    .cast_valid_i_7_23                              (cast_valid_pe_2_nw[7][23]),
    .cast_ready_o_7_23                              (cast_ready_nw_2_pe[7][23]),
    .merge_data_i_7_23                              (merge_data_pe_2_nw[7][23]),
    .merge_valid_i_7_23                             (merge_valid_pe_2_nw[7][23]),
    .merge_ready_o_7_23                             (merge_ready_nw_2_pe[7][23]),
    .gather_data_i_7_23                             (gather_data_pe_2_nw[7][23]),
    .gather_valid_i_7_23                            (gather_valid_pe_2_nw[7][23]),
    .gather_ready_o_7_23                            (gather_ready_nw_2_pe[7][23]),

    .cast_data_o_7_23                               (cast_data_nw_2_pe[7][23]),
    .cast_valid_o_7_23                              (cast_valid_nw_2_pe[7][23]),
    .cast_ready_i_7_23                              (cast_ready_pe_2_nw[7][23]),
    .merge_data_o_7_23                              (merge_data_nw_2_pe[7][23]),
    .merge_valid_o_7_23                             (merge_valid_nw_2_pe[7][23]),
    .merge_ready_i_7_23                             (merge_ready_pe_2_nw[7][23]),
    .gather_data_o_7_23                             (gather_data_nw_2_pe[7][23]),
    .gather_valid_o_7_23                            (gather_valid_nw_2_pe[7][23]),
    .gather_ready_i_7_23                            (gather_ready_pe_2_nw[7][23]),
    .cast_data_i_7_24                               (cast_data_pe_2_nw[7][24]),
    .cast_valid_i_7_24                              (cast_valid_pe_2_nw[7][24]),
    .cast_ready_o_7_24                              (cast_ready_nw_2_pe[7][24]),
    .merge_data_i_7_24                              (merge_data_pe_2_nw[7][24]),
    .merge_valid_i_7_24                             (merge_valid_pe_2_nw[7][24]),
    .merge_ready_o_7_24                             (merge_ready_nw_2_pe[7][24]),
    .gather_data_i_7_24                             (gather_data_pe_2_nw[7][24]),
    .gather_valid_i_7_24                            (gather_valid_pe_2_nw[7][24]),
    .gather_ready_o_7_24                            (gather_ready_nw_2_pe[7][24]),

    .cast_data_o_7_24                               (cast_data_nw_2_pe[7][24]),
    .cast_valid_o_7_24                              (cast_valid_nw_2_pe[7][24]),
    .cast_ready_i_7_24                              (cast_ready_pe_2_nw[7][24]),
    .merge_data_o_7_24                              (merge_data_nw_2_pe[7][24]),
    .merge_valid_o_7_24                             (merge_valid_nw_2_pe[7][24]),
    .merge_ready_i_7_24                             (merge_ready_pe_2_nw[7][24]),
    .gather_data_o_7_24                             (gather_data_nw_2_pe[7][24]),
    .gather_valid_o_7_24                            (gather_valid_nw_2_pe[7][24]),
    .gather_ready_i_7_24                            (gather_ready_pe_2_nw[7][24]),
    .cast_data_i_8_0                               (cast_data_pe_2_nw[8][0]),
    .cast_valid_i_8_0                              (cast_valid_pe_2_nw[8][0]),
    .cast_ready_o_8_0                              (cast_ready_nw_2_pe[8][0]),
    .merge_data_i_8_0                              (merge_data_pe_2_nw[8][0]),
    .merge_valid_i_8_0                             (merge_valid_pe_2_nw[8][0]),
    .merge_ready_o_8_0                             (merge_ready_nw_2_pe[8][0]),
    .gather_data_i_8_0                             (gather_data_pe_2_nw[8][0]),
    .gather_valid_i_8_0                            (gather_valid_pe_2_nw[8][0]),
    .gather_ready_o_8_0                            (gather_ready_nw_2_pe[8][0]),

    .cast_data_o_8_0                               (cast_data_nw_2_pe[8][0]),
    .cast_valid_o_8_0                              (cast_valid_nw_2_pe[8][0]),
    .cast_ready_i_8_0                              (cast_ready_pe_2_nw[8][0]),
    .merge_data_o_8_0                              (merge_data_nw_2_pe[8][0]),
    .merge_valid_o_8_0                             (merge_valid_nw_2_pe[8][0]),
    .merge_ready_i_8_0                             (merge_ready_pe_2_nw[8][0]),
    .gather_data_o_8_0                             (gather_data_nw_2_pe[8][0]),
    .gather_valid_o_8_0                            (gather_valid_nw_2_pe[8][0]),
    .gather_ready_i_8_0                            (gather_ready_pe_2_nw[8][0]),
    .cast_data_i_8_1                               (cast_data_pe_2_nw[8][1]),
    .cast_valid_i_8_1                              (cast_valid_pe_2_nw[8][1]),
    .cast_ready_o_8_1                              (cast_ready_nw_2_pe[8][1]),
    .merge_data_i_8_1                              (merge_data_pe_2_nw[8][1]),
    .merge_valid_i_8_1                             (merge_valid_pe_2_nw[8][1]),
    .merge_ready_o_8_1                             (merge_ready_nw_2_pe[8][1]),
    .gather_data_i_8_1                             (gather_data_pe_2_nw[8][1]),
    .gather_valid_i_8_1                            (gather_valid_pe_2_nw[8][1]),
    .gather_ready_o_8_1                            (gather_ready_nw_2_pe[8][1]),

    .cast_data_o_8_1                               (cast_data_nw_2_pe[8][1]),
    .cast_valid_o_8_1                              (cast_valid_nw_2_pe[8][1]),
    .cast_ready_i_8_1                              (cast_ready_pe_2_nw[8][1]),
    .merge_data_o_8_1                              (merge_data_nw_2_pe[8][1]),
    .merge_valid_o_8_1                             (merge_valid_nw_2_pe[8][1]),
    .merge_ready_i_8_1                             (merge_ready_pe_2_nw[8][1]),
    .gather_data_o_8_1                             (gather_data_nw_2_pe[8][1]),
    .gather_valid_o_8_1                            (gather_valid_nw_2_pe[8][1]),
    .gather_ready_i_8_1                            (gather_ready_pe_2_nw[8][1]),
    .cast_data_i_8_2                               (cast_data_pe_2_nw[8][2]),
    .cast_valid_i_8_2                              (cast_valid_pe_2_nw[8][2]),
    .cast_ready_o_8_2                              (cast_ready_nw_2_pe[8][2]),
    .merge_data_i_8_2                              (merge_data_pe_2_nw[8][2]),
    .merge_valid_i_8_2                             (merge_valid_pe_2_nw[8][2]),
    .merge_ready_o_8_2                             (merge_ready_nw_2_pe[8][2]),
    .gather_data_i_8_2                             (gather_data_pe_2_nw[8][2]),
    .gather_valid_i_8_2                            (gather_valid_pe_2_nw[8][2]),
    .gather_ready_o_8_2                            (gather_ready_nw_2_pe[8][2]),

    .cast_data_o_8_2                               (cast_data_nw_2_pe[8][2]),
    .cast_valid_o_8_2                              (cast_valid_nw_2_pe[8][2]),
    .cast_ready_i_8_2                              (cast_ready_pe_2_nw[8][2]),
    .merge_data_o_8_2                              (merge_data_nw_2_pe[8][2]),
    .merge_valid_o_8_2                             (merge_valid_nw_2_pe[8][2]),
    .merge_ready_i_8_2                             (merge_ready_pe_2_nw[8][2]),
    .gather_data_o_8_2                             (gather_data_nw_2_pe[8][2]),
    .gather_valid_o_8_2                            (gather_valid_nw_2_pe[8][2]),
    .gather_ready_i_8_2                            (gather_ready_pe_2_nw[8][2]),
    .cast_data_i_8_3                               (cast_data_pe_2_nw[8][3]),
    .cast_valid_i_8_3                              (cast_valid_pe_2_nw[8][3]),
    .cast_ready_o_8_3                              (cast_ready_nw_2_pe[8][3]),
    .merge_data_i_8_3                              (merge_data_pe_2_nw[8][3]),
    .merge_valid_i_8_3                             (merge_valid_pe_2_nw[8][3]),
    .merge_ready_o_8_3                             (merge_ready_nw_2_pe[8][3]),
    .gather_data_i_8_3                             (gather_data_pe_2_nw[8][3]),
    .gather_valid_i_8_3                            (gather_valid_pe_2_nw[8][3]),
    .gather_ready_o_8_3                            (gather_ready_nw_2_pe[8][3]),

    .cast_data_o_8_3                               (cast_data_nw_2_pe[8][3]),
    .cast_valid_o_8_3                              (cast_valid_nw_2_pe[8][3]),
    .cast_ready_i_8_3                              (cast_ready_pe_2_nw[8][3]),
    .merge_data_o_8_3                              (merge_data_nw_2_pe[8][3]),
    .merge_valid_o_8_3                             (merge_valid_nw_2_pe[8][3]),
    .merge_ready_i_8_3                             (merge_ready_pe_2_nw[8][3]),
    .gather_data_o_8_3                             (gather_data_nw_2_pe[8][3]),
    .gather_valid_o_8_3                            (gather_valid_nw_2_pe[8][3]),
    .gather_ready_i_8_3                            (gather_ready_pe_2_nw[8][3]),
    .cast_data_i_8_4                               (cast_data_pe_2_nw[8][4]),
    .cast_valid_i_8_4                              (cast_valid_pe_2_nw[8][4]),
    .cast_ready_o_8_4                              (cast_ready_nw_2_pe[8][4]),
    .merge_data_i_8_4                              (merge_data_pe_2_nw[8][4]),
    .merge_valid_i_8_4                             (merge_valid_pe_2_nw[8][4]),
    .merge_ready_o_8_4                             (merge_ready_nw_2_pe[8][4]),
    .gather_data_i_8_4                             (gather_data_pe_2_nw[8][4]),
    .gather_valid_i_8_4                            (gather_valid_pe_2_nw[8][4]),
    .gather_ready_o_8_4                            (gather_ready_nw_2_pe[8][4]),

    .cast_data_o_8_4                               (cast_data_nw_2_pe[8][4]),
    .cast_valid_o_8_4                              (cast_valid_nw_2_pe[8][4]),
    .cast_ready_i_8_4                              (cast_ready_pe_2_nw[8][4]),
    .merge_data_o_8_4                              (merge_data_nw_2_pe[8][4]),
    .merge_valid_o_8_4                             (merge_valid_nw_2_pe[8][4]),
    .merge_ready_i_8_4                             (merge_ready_pe_2_nw[8][4]),
    .gather_data_o_8_4                             (gather_data_nw_2_pe[8][4]),
    .gather_valid_o_8_4                            (gather_valid_nw_2_pe[8][4]),
    .gather_ready_i_8_4                            (gather_ready_pe_2_nw[8][4]),
    .cast_data_i_8_5                               (cast_data_pe_2_nw[8][5]),
    .cast_valid_i_8_5                              (cast_valid_pe_2_nw[8][5]),
    .cast_ready_o_8_5                              (cast_ready_nw_2_pe[8][5]),
    .merge_data_i_8_5                              (merge_data_pe_2_nw[8][5]),
    .merge_valid_i_8_5                             (merge_valid_pe_2_nw[8][5]),
    .merge_ready_o_8_5                             (merge_ready_nw_2_pe[8][5]),
    .gather_data_i_8_5                             (gather_data_pe_2_nw[8][5]),
    .gather_valid_i_8_5                            (gather_valid_pe_2_nw[8][5]),
    .gather_ready_o_8_5                            (gather_ready_nw_2_pe[8][5]),

    .cast_data_o_8_5                               (cast_data_nw_2_pe[8][5]),
    .cast_valid_o_8_5                              (cast_valid_nw_2_pe[8][5]),
    .cast_ready_i_8_5                              (cast_ready_pe_2_nw[8][5]),
    .merge_data_o_8_5                              (merge_data_nw_2_pe[8][5]),
    .merge_valid_o_8_5                             (merge_valid_nw_2_pe[8][5]),
    .merge_ready_i_8_5                             (merge_ready_pe_2_nw[8][5]),
    .gather_data_o_8_5                             (gather_data_nw_2_pe[8][5]),
    .gather_valid_o_8_5                            (gather_valid_nw_2_pe[8][5]),
    .gather_ready_i_8_5                            (gather_ready_pe_2_nw[8][5]),
    .cast_data_i_8_6                               (cast_data_pe_2_nw[8][6]),
    .cast_valid_i_8_6                              (cast_valid_pe_2_nw[8][6]),
    .cast_ready_o_8_6                              (cast_ready_nw_2_pe[8][6]),
    .merge_data_i_8_6                              (merge_data_pe_2_nw[8][6]),
    .merge_valid_i_8_6                             (merge_valid_pe_2_nw[8][6]),
    .merge_ready_o_8_6                             (merge_ready_nw_2_pe[8][6]),
    .gather_data_i_8_6                             (gather_data_pe_2_nw[8][6]),
    .gather_valid_i_8_6                            (gather_valid_pe_2_nw[8][6]),
    .gather_ready_o_8_6                            (gather_ready_nw_2_pe[8][6]),

    .cast_data_o_8_6                               (cast_data_nw_2_pe[8][6]),
    .cast_valid_o_8_6                              (cast_valid_nw_2_pe[8][6]),
    .cast_ready_i_8_6                              (cast_ready_pe_2_nw[8][6]),
    .merge_data_o_8_6                              (merge_data_nw_2_pe[8][6]),
    .merge_valid_o_8_6                             (merge_valid_nw_2_pe[8][6]),
    .merge_ready_i_8_6                             (merge_ready_pe_2_nw[8][6]),
    .gather_data_o_8_6                             (gather_data_nw_2_pe[8][6]),
    .gather_valid_o_8_6                            (gather_valid_nw_2_pe[8][6]),
    .gather_ready_i_8_6                            (gather_ready_pe_2_nw[8][6]),
    .cast_data_i_8_7                               (cast_data_pe_2_nw[8][7]),
    .cast_valid_i_8_7                              (cast_valid_pe_2_nw[8][7]),
    .cast_ready_o_8_7                              (cast_ready_nw_2_pe[8][7]),
    .merge_data_i_8_7                              (merge_data_pe_2_nw[8][7]),
    .merge_valid_i_8_7                             (merge_valid_pe_2_nw[8][7]),
    .merge_ready_o_8_7                             (merge_ready_nw_2_pe[8][7]),
    .gather_data_i_8_7                             (gather_data_pe_2_nw[8][7]),
    .gather_valid_i_8_7                            (gather_valid_pe_2_nw[8][7]),
    .gather_ready_o_8_7                            (gather_ready_nw_2_pe[8][7]),

    .cast_data_o_8_7                               (cast_data_nw_2_pe[8][7]),
    .cast_valid_o_8_7                              (cast_valid_nw_2_pe[8][7]),
    .cast_ready_i_8_7                              (cast_ready_pe_2_nw[8][7]),
    .merge_data_o_8_7                              (merge_data_nw_2_pe[8][7]),
    .merge_valid_o_8_7                             (merge_valid_nw_2_pe[8][7]),
    .merge_ready_i_8_7                             (merge_ready_pe_2_nw[8][7]),
    .gather_data_o_8_7                             (gather_data_nw_2_pe[8][7]),
    .gather_valid_o_8_7                            (gather_valid_nw_2_pe[8][7]),
    .gather_ready_i_8_7                            (gather_ready_pe_2_nw[8][7]),
    .cast_data_i_8_8                               (cast_data_pe_2_nw[8][8]),
    .cast_valid_i_8_8                              (cast_valid_pe_2_nw[8][8]),
    .cast_ready_o_8_8                              (cast_ready_nw_2_pe[8][8]),
    .merge_data_i_8_8                              (merge_data_pe_2_nw[8][8]),
    .merge_valid_i_8_8                             (merge_valid_pe_2_nw[8][8]),
    .merge_ready_o_8_8                             (merge_ready_nw_2_pe[8][8]),
    .gather_data_i_8_8                             (gather_data_pe_2_nw[8][8]),
    .gather_valid_i_8_8                            (gather_valid_pe_2_nw[8][8]),
    .gather_ready_o_8_8                            (gather_ready_nw_2_pe[8][8]),

    .cast_data_o_8_8                               (cast_data_nw_2_pe[8][8]),
    .cast_valid_o_8_8                              (cast_valid_nw_2_pe[8][8]),
    .cast_ready_i_8_8                              (cast_ready_pe_2_nw[8][8]),
    .merge_data_o_8_8                              (merge_data_nw_2_pe[8][8]),
    .merge_valid_o_8_8                             (merge_valid_nw_2_pe[8][8]),
    .merge_ready_i_8_8                             (merge_ready_pe_2_nw[8][8]),
    .gather_data_o_8_8                             (gather_data_nw_2_pe[8][8]),
    .gather_valid_o_8_8                            (gather_valid_nw_2_pe[8][8]),
    .gather_ready_i_8_8                            (gather_ready_pe_2_nw[8][8]),
    .cast_data_i_8_9                               (cast_data_pe_2_nw[8][9]),
    .cast_valid_i_8_9                              (cast_valid_pe_2_nw[8][9]),
    .cast_ready_o_8_9                              (cast_ready_nw_2_pe[8][9]),
    .merge_data_i_8_9                              (merge_data_pe_2_nw[8][9]),
    .merge_valid_i_8_9                             (merge_valid_pe_2_nw[8][9]),
    .merge_ready_o_8_9                             (merge_ready_nw_2_pe[8][9]),
    .gather_data_i_8_9                             (gather_data_pe_2_nw[8][9]),
    .gather_valid_i_8_9                            (gather_valid_pe_2_nw[8][9]),
    .gather_ready_o_8_9                            (gather_ready_nw_2_pe[8][9]),

    .cast_data_o_8_9                               (cast_data_nw_2_pe[8][9]),
    .cast_valid_o_8_9                              (cast_valid_nw_2_pe[8][9]),
    .cast_ready_i_8_9                              (cast_ready_pe_2_nw[8][9]),
    .merge_data_o_8_9                              (merge_data_nw_2_pe[8][9]),
    .merge_valid_o_8_9                             (merge_valid_nw_2_pe[8][9]),
    .merge_ready_i_8_9                             (merge_ready_pe_2_nw[8][9]),
    .gather_data_o_8_9                             (gather_data_nw_2_pe[8][9]),
    .gather_valid_o_8_9                            (gather_valid_nw_2_pe[8][9]),
    .gather_ready_i_8_9                            (gather_ready_pe_2_nw[8][9]),
    .cast_data_i_8_10                               (cast_data_pe_2_nw[8][10]),
    .cast_valid_i_8_10                              (cast_valid_pe_2_nw[8][10]),
    .cast_ready_o_8_10                              (cast_ready_nw_2_pe[8][10]),
    .merge_data_i_8_10                              (merge_data_pe_2_nw[8][10]),
    .merge_valid_i_8_10                             (merge_valid_pe_2_nw[8][10]),
    .merge_ready_o_8_10                             (merge_ready_nw_2_pe[8][10]),
    .gather_data_i_8_10                             (gather_data_pe_2_nw[8][10]),
    .gather_valid_i_8_10                            (gather_valid_pe_2_nw[8][10]),
    .gather_ready_o_8_10                            (gather_ready_nw_2_pe[8][10]),

    .cast_data_o_8_10                               (cast_data_nw_2_pe[8][10]),
    .cast_valid_o_8_10                              (cast_valid_nw_2_pe[8][10]),
    .cast_ready_i_8_10                              (cast_ready_pe_2_nw[8][10]),
    .merge_data_o_8_10                              (merge_data_nw_2_pe[8][10]),
    .merge_valid_o_8_10                             (merge_valid_nw_2_pe[8][10]),
    .merge_ready_i_8_10                             (merge_ready_pe_2_nw[8][10]),
    .gather_data_o_8_10                             (gather_data_nw_2_pe[8][10]),
    .gather_valid_o_8_10                            (gather_valid_nw_2_pe[8][10]),
    .gather_ready_i_8_10                            (gather_ready_pe_2_nw[8][10]),
    .cast_data_i_8_11                               (cast_data_pe_2_nw[8][11]),
    .cast_valid_i_8_11                              (cast_valid_pe_2_nw[8][11]),
    .cast_ready_o_8_11                              (cast_ready_nw_2_pe[8][11]),
    .merge_data_i_8_11                              (merge_data_pe_2_nw[8][11]),
    .merge_valid_i_8_11                             (merge_valid_pe_2_nw[8][11]),
    .merge_ready_o_8_11                             (merge_ready_nw_2_pe[8][11]),
    .gather_data_i_8_11                             (gather_data_pe_2_nw[8][11]),
    .gather_valid_i_8_11                            (gather_valid_pe_2_nw[8][11]),
    .gather_ready_o_8_11                            (gather_ready_nw_2_pe[8][11]),

    .cast_data_o_8_11                               (cast_data_nw_2_pe[8][11]),
    .cast_valid_o_8_11                              (cast_valid_nw_2_pe[8][11]),
    .cast_ready_i_8_11                              (cast_ready_pe_2_nw[8][11]),
    .merge_data_o_8_11                              (merge_data_nw_2_pe[8][11]),
    .merge_valid_o_8_11                             (merge_valid_nw_2_pe[8][11]),
    .merge_ready_i_8_11                             (merge_ready_pe_2_nw[8][11]),
    .gather_data_o_8_11                             (gather_data_nw_2_pe[8][11]),
    .gather_valid_o_8_11                            (gather_valid_nw_2_pe[8][11]),
    .gather_ready_i_8_11                            (gather_ready_pe_2_nw[8][11]),
    .cast_data_i_8_12                               (cast_data_pe_2_nw[8][12]),
    .cast_valid_i_8_12                              (cast_valid_pe_2_nw[8][12]),
    .cast_ready_o_8_12                              (cast_ready_nw_2_pe[8][12]),
    .merge_data_i_8_12                              (merge_data_pe_2_nw[8][12]),
    .merge_valid_i_8_12                             (merge_valid_pe_2_nw[8][12]),
    .merge_ready_o_8_12                             (merge_ready_nw_2_pe[8][12]),
    .gather_data_i_8_12                             (gather_data_pe_2_nw[8][12]),
    .gather_valid_i_8_12                            (gather_valid_pe_2_nw[8][12]),
    .gather_ready_o_8_12                            (gather_ready_nw_2_pe[8][12]),

    .cast_data_o_8_12                               (cast_data_nw_2_pe[8][12]),
    .cast_valid_o_8_12                              (cast_valid_nw_2_pe[8][12]),
    .cast_ready_i_8_12                              (cast_ready_pe_2_nw[8][12]),
    .merge_data_o_8_12                              (merge_data_nw_2_pe[8][12]),
    .merge_valid_o_8_12                             (merge_valid_nw_2_pe[8][12]),
    .merge_ready_i_8_12                             (merge_ready_pe_2_nw[8][12]),
    .gather_data_o_8_12                             (gather_data_nw_2_pe[8][12]),
    .gather_valid_o_8_12                            (gather_valid_nw_2_pe[8][12]),
    .gather_ready_i_8_12                            (gather_ready_pe_2_nw[8][12]),
    .cast_data_i_8_13                               (cast_data_pe_2_nw[8][13]),
    .cast_valid_i_8_13                              (cast_valid_pe_2_nw[8][13]),
    .cast_ready_o_8_13                              (cast_ready_nw_2_pe[8][13]),
    .merge_data_i_8_13                              (merge_data_pe_2_nw[8][13]),
    .merge_valid_i_8_13                             (merge_valid_pe_2_nw[8][13]),
    .merge_ready_o_8_13                             (merge_ready_nw_2_pe[8][13]),
    .gather_data_i_8_13                             (gather_data_pe_2_nw[8][13]),
    .gather_valid_i_8_13                            (gather_valid_pe_2_nw[8][13]),
    .gather_ready_o_8_13                            (gather_ready_nw_2_pe[8][13]),

    .cast_data_o_8_13                               (cast_data_nw_2_pe[8][13]),
    .cast_valid_o_8_13                              (cast_valid_nw_2_pe[8][13]),
    .cast_ready_i_8_13                              (cast_ready_pe_2_nw[8][13]),
    .merge_data_o_8_13                              (merge_data_nw_2_pe[8][13]),
    .merge_valid_o_8_13                             (merge_valid_nw_2_pe[8][13]),
    .merge_ready_i_8_13                             (merge_ready_pe_2_nw[8][13]),
    .gather_data_o_8_13                             (gather_data_nw_2_pe[8][13]),
    .gather_valid_o_8_13                            (gather_valid_nw_2_pe[8][13]),
    .gather_ready_i_8_13                            (gather_ready_pe_2_nw[8][13]),
    .cast_data_i_8_14                               (cast_data_pe_2_nw[8][14]),
    .cast_valid_i_8_14                              (cast_valid_pe_2_nw[8][14]),
    .cast_ready_o_8_14                              (cast_ready_nw_2_pe[8][14]),
    .merge_data_i_8_14                              (merge_data_pe_2_nw[8][14]),
    .merge_valid_i_8_14                             (merge_valid_pe_2_nw[8][14]),
    .merge_ready_o_8_14                             (merge_ready_nw_2_pe[8][14]),
    .gather_data_i_8_14                             (gather_data_pe_2_nw[8][14]),
    .gather_valid_i_8_14                            (gather_valid_pe_2_nw[8][14]),
    .gather_ready_o_8_14                            (gather_ready_nw_2_pe[8][14]),

    .cast_data_o_8_14                               (cast_data_nw_2_pe[8][14]),
    .cast_valid_o_8_14                              (cast_valid_nw_2_pe[8][14]),
    .cast_ready_i_8_14                              (cast_ready_pe_2_nw[8][14]),
    .merge_data_o_8_14                              (merge_data_nw_2_pe[8][14]),
    .merge_valid_o_8_14                             (merge_valid_nw_2_pe[8][14]),
    .merge_ready_i_8_14                             (merge_ready_pe_2_nw[8][14]),
    .gather_data_o_8_14                             (gather_data_nw_2_pe[8][14]),
    .gather_valid_o_8_14                            (gather_valid_nw_2_pe[8][14]),
    .gather_ready_i_8_14                            (gather_ready_pe_2_nw[8][14]),
    .cast_data_i_8_15                               (cast_data_pe_2_nw[8][15]),
    .cast_valid_i_8_15                              (cast_valid_pe_2_nw[8][15]),
    .cast_ready_o_8_15                              (cast_ready_nw_2_pe[8][15]),
    .merge_data_i_8_15                              (merge_data_pe_2_nw[8][15]),
    .merge_valid_i_8_15                             (merge_valid_pe_2_nw[8][15]),
    .merge_ready_o_8_15                             (merge_ready_nw_2_pe[8][15]),
    .gather_data_i_8_15                             (gather_data_pe_2_nw[8][15]),
    .gather_valid_i_8_15                            (gather_valid_pe_2_nw[8][15]),
    .gather_ready_o_8_15                            (gather_ready_nw_2_pe[8][15]),

    .cast_data_o_8_15                               (cast_data_nw_2_pe[8][15]),
    .cast_valid_o_8_15                              (cast_valid_nw_2_pe[8][15]),
    .cast_ready_i_8_15                              (cast_ready_pe_2_nw[8][15]),
    .merge_data_o_8_15                              (merge_data_nw_2_pe[8][15]),
    .merge_valid_o_8_15                             (merge_valid_nw_2_pe[8][15]),
    .merge_ready_i_8_15                             (merge_ready_pe_2_nw[8][15]),
    .gather_data_o_8_15                             (gather_data_nw_2_pe[8][15]),
    .gather_valid_o_8_15                            (gather_valid_nw_2_pe[8][15]),
    .gather_ready_i_8_15                            (gather_ready_pe_2_nw[8][15]),
    .cast_data_i_8_16                               (cast_data_pe_2_nw[8][16]),
    .cast_valid_i_8_16                              (cast_valid_pe_2_nw[8][16]),
    .cast_ready_o_8_16                              (cast_ready_nw_2_pe[8][16]),
    .merge_data_i_8_16                              (merge_data_pe_2_nw[8][16]),
    .merge_valid_i_8_16                             (merge_valid_pe_2_nw[8][16]),
    .merge_ready_o_8_16                             (merge_ready_nw_2_pe[8][16]),
    .gather_data_i_8_16                             (gather_data_pe_2_nw[8][16]),
    .gather_valid_i_8_16                            (gather_valid_pe_2_nw[8][16]),
    .gather_ready_o_8_16                            (gather_ready_nw_2_pe[8][16]),

    .cast_data_o_8_16                               (cast_data_nw_2_pe[8][16]),
    .cast_valid_o_8_16                              (cast_valid_nw_2_pe[8][16]),
    .cast_ready_i_8_16                              (cast_ready_pe_2_nw[8][16]),
    .merge_data_o_8_16                              (merge_data_nw_2_pe[8][16]),
    .merge_valid_o_8_16                             (merge_valid_nw_2_pe[8][16]),
    .merge_ready_i_8_16                             (merge_ready_pe_2_nw[8][16]),
    .gather_data_o_8_16                             (gather_data_nw_2_pe[8][16]),
    .gather_valid_o_8_16                            (gather_valid_nw_2_pe[8][16]),
    .gather_ready_i_8_16                            (gather_ready_pe_2_nw[8][16]),
    .cast_data_i_8_17                               (cast_data_pe_2_nw[8][17]),
    .cast_valid_i_8_17                              (cast_valid_pe_2_nw[8][17]),
    .cast_ready_o_8_17                              (cast_ready_nw_2_pe[8][17]),
    .merge_data_i_8_17                              (merge_data_pe_2_nw[8][17]),
    .merge_valid_i_8_17                             (merge_valid_pe_2_nw[8][17]),
    .merge_ready_o_8_17                             (merge_ready_nw_2_pe[8][17]),
    .gather_data_i_8_17                             (gather_data_pe_2_nw[8][17]),
    .gather_valid_i_8_17                            (gather_valid_pe_2_nw[8][17]),
    .gather_ready_o_8_17                            (gather_ready_nw_2_pe[8][17]),

    .cast_data_o_8_17                               (cast_data_nw_2_pe[8][17]),
    .cast_valid_o_8_17                              (cast_valid_nw_2_pe[8][17]),
    .cast_ready_i_8_17                              (cast_ready_pe_2_nw[8][17]),
    .merge_data_o_8_17                              (merge_data_nw_2_pe[8][17]),
    .merge_valid_o_8_17                             (merge_valid_nw_2_pe[8][17]),
    .merge_ready_i_8_17                             (merge_ready_pe_2_nw[8][17]),
    .gather_data_o_8_17                             (gather_data_nw_2_pe[8][17]),
    .gather_valid_o_8_17                            (gather_valid_nw_2_pe[8][17]),
    .gather_ready_i_8_17                            (gather_ready_pe_2_nw[8][17]),
    .cast_data_i_8_18                               (cast_data_pe_2_nw[8][18]),
    .cast_valid_i_8_18                              (cast_valid_pe_2_nw[8][18]),
    .cast_ready_o_8_18                              (cast_ready_nw_2_pe[8][18]),
    .merge_data_i_8_18                              (merge_data_pe_2_nw[8][18]),
    .merge_valid_i_8_18                             (merge_valid_pe_2_nw[8][18]),
    .merge_ready_o_8_18                             (merge_ready_nw_2_pe[8][18]),
    .gather_data_i_8_18                             (gather_data_pe_2_nw[8][18]),
    .gather_valid_i_8_18                            (gather_valid_pe_2_nw[8][18]),
    .gather_ready_o_8_18                            (gather_ready_nw_2_pe[8][18]),

    .cast_data_o_8_18                               (cast_data_nw_2_pe[8][18]),
    .cast_valid_o_8_18                              (cast_valid_nw_2_pe[8][18]),
    .cast_ready_i_8_18                              (cast_ready_pe_2_nw[8][18]),
    .merge_data_o_8_18                              (merge_data_nw_2_pe[8][18]),
    .merge_valid_o_8_18                             (merge_valid_nw_2_pe[8][18]),
    .merge_ready_i_8_18                             (merge_ready_pe_2_nw[8][18]),
    .gather_data_o_8_18                             (gather_data_nw_2_pe[8][18]),
    .gather_valid_o_8_18                            (gather_valid_nw_2_pe[8][18]),
    .gather_ready_i_8_18                            (gather_ready_pe_2_nw[8][18]),
    .cast_data_i_8_19                               (cast_data_pe_2_nw[8][19]),
    .cast_valid_i_8_19                              (cast_valid_pe_2_nw[8][19]),
    .cast_ready_o_8_19                              (cast_ready_nw_2_pe[8][19]),
    .merge_data_i_8_19                              (merge_data_pe_2_nw[8][19]),
    .merge_valid_i_8_19                             (merge_valid_pe_2_nw[8][19]),
    .merge_ready_o_8_19                             (merge_ready_nw_2_pe[8][19]),
    .gather_data_i_8_19                             (gather_data_pe_2_nw[8][19]),
    .gather_valid_i_8_19                            (gather_valid_pe_2_nw[8][19]),
    .gather_ready_o_8_19                            (gather_ready_nw_2_pe[8][19]),

    .cast_data_o_8_19                               (cast_data_nw_2_pe[8][19]),
    .cast_valid_o_8_19                              (cast_valid_nw_2_pe[8][19]),
    .cast_ready_i_8_19                              (cast_ready_pe_2_nw[8][19]),
    .merge_data_o_8_19                              (merge_data_nw_2_pe[8][19]),
    .merge_valid_o_8_19                             (merge_valid_nw_2_pe[8][19]),
    .merge_ready_i_8_19                             (merge_ready_pe_2_nw[8][19]),
    .gather_data_o_8_19                             (gather_data_nw_2_pe[8][19]),
    .gather_valid_o_8_19                            (gather_valid_nw_2_pe[8][19]),
    .gather_ready_i_8_19                            (gather_ready_pe_2_nw[8][19]),
    .cast_data_i_8_20                               (cast_data_pe_2_nw[8][20]),
    .cast_valid_i_8_20                              (cast_valid_pe_2_nw[8][20]),
    .cast_ready_o_8_20                              (cast_ready_nw_2_pe[8][20]),
    .merge_data_i_8_20                              (merge_data_pe_2_nw[8][20]),
    .merge_valid_i_8_20                             (merge_valid_pe_2_nw[8][20]),
    .merge_ready_o_8_20                             (merge_ready_nw_2_pe[8][20]),
    .gather_data_i_8_20                             (gather_data_pe_2_nw[8][20]),
    .gather_valid_i_8_20                            (gather_valid_pe_2_nw[8][20]),
    .gather_ready_o_8_20                            (gather_ready_nw_2_pe[8][20]),

    .cast_data_o_8_20                               (cast_data_nw_2_pe[8][20]),
    .cast_valid_o_8_20                              (cast_valid_nw_2_pe[8][20]),
    .cast_ready_i_8_20                              (cast_ready_pe_2_nw[8][20]),
    .merge_data_o_8_20                              (merge_data_nw_2_pe[8][20]),
    .merge_valid_o_8_20                             (merge_valid_nw_2_pe[8][20]),
    .merge_ready_i_8_20                             (merge_ready_pe_2_nw[8][20]),
    .gather_data_o_8_20                             (gather_data_nw_2_pe[8][20]),
    .gather_valid_o_8_20                            (gather_valid_nw_2_pe[8][20]),
    .gather_ready_i_8_20                            (gather_ready_pe_2_nw[8][20]),
    .cast_data_i_8_21                               (cast_data_pe_2_nw[8][21]),
    .cast_valid_i_8_21                              (cast_valid_pe_2_nw[8][21]),
    .cast_ready_o_8_21                              (cast_ready_nw_2_pe[8][21]),
    .merge_data_i_8_21                              (merge_data_pe_2_nw[8][21]),
    .merge_valid_i_8_21                             (merge_valid_pe_2_nw[8][21]),
    .merge_ready_o_8_21                             (merge_ready_nw_2_pe[8][21]),
    .gather_data_i_8_21                             (gather_data_pe_2_nw[8][21]),
    .gather_valid_i_8_21                            (gather_valid_pe_2_nw[8][21]),
    .gather_ready_o_8_21                            (gather_ready_nw_2_pe[8][21]),

    .cast_data_o_8_21                               (cast_data_nw_2_pe[8][21]),
    .cast_valid_o_8_21                              (cast_valid_nw_2_pe[8][21]),
    .cast_ready_i_8_21                              (cast_ready_pe_2_nw[8][21]),
    .merge_data_o_8_21                              (merge_data_nw_2_pe[8][21]),
    .merge_valid_o_8_21                             (merge_valid_nw_2_pe[8][21]),
    .merge_ready_i_8_21                             (merge_ready_pe_2_nw[8][21]),
    .gather_data_o_8_21                             (gather_data_nw_2_pe[8][21]),
    .gather_valid_o_8_21                            (gather_valid_nw_2_pe[8][21]),
    .gather_ready_i_8_21                            (gather_ready_pe_2_nw[8][21]),
    .cast_data_i_8_22                               (cast_data_pe_2_nw[8][22]),
    .cast_valid_i_8_22                              (cast_valid_pe_2_nw[8][22]),
    .cast_ready_o_8_22                              (cast_ready_nw_2_pe[8][22]),
    .merge_data_i_8_22                              (merge_data_pe_2_nw[8][22]),
    .merge_valid_i_8_22                             (merge_valid_pe_2_nw[8][22]),
    .merge_ready_o_8_22                             (merge_ready_nw_2_pe[8][22]),
    .gather_data_i_8_22                             (gather_data_pe_2_nw[8][22]),
    .gather_valid_i_8_22                            (gather_valid_pe_2_nw[8][22]),
    .gather_ready_o_8_22                            (gather_ready_nw_2_pe[8][22]),

    .cast_data_o_8_22                               (cast_data_nw_2_pe[8][22]),
    .cast_valid_o_8_22                              (cast_valid_nw_2_pe[8][22]),
    .cast_ready_i_8_22                              (cast_ready_pe_2_nw[8][22]),
    .merge_data_o_8_22                              (merge_data_nw_2_pe[8][22]),
    .merge_valid_o_8_22                             (merge_valid_nw_2_pe[8][22]),
    .merge_ready_i_8_22                             (merge_ready_pe_2_nw[8][22]),
    .gather_data_o_8_22                             (gather_data_nw_2_pe[8][22]),
    .gather_valid_o_8_22                            (gather_valid_nw_2_pe[8][22]),
    .gather_ready_i_8_22                            (gather_ready_pe_2_nw[8][22]),
    .cast_data_i_8_23                               (cast_data_pe_2_nw[8][23]),
    .cast_valid_i_8_23                              (cast_valid_pe_2_nw[8][23]),
    .cast_ready_o_8_23                              (cast_ready_nw_2_pe[8][23]),
    .merge_data_i_8_23                              (merge_data_pe_2_nw[8][23]),
    .merge_valid_i_8_23                             (merge_valid_pe_2_nw[8][23]),
    .merge_ready_o_8_23                             (merge_ready_nw_2_pe[8][23]),
    .gather_data_i_8_23                             (gather_data_pe_2_nw[8][23]),
    .gather_valid_i_8_23                            (gather_valid_pe_2_nw[8][23]),
    .gather_ready_o_8_23                            (gather_ready_nw_2_pe[8][23]),

    .cast_data_o_8_23                               (cast_data_nw_2_pe[8][23]),
    .cast_valid_o_8_23                              (cast_valid_nw_2_pe[8][23]),
    .cast_ready_i_8_23                              (cast_ready_pe_2_nw[8][23]),
    .merge_data_o_8_23                              (merge_data_nw_2_pe[8][23]),
    .merge_valid_o_8_23                             (merge_valid_nw_2_pe[8][23]),
    .merge_ready_i_8_23                             (merge_ready_pe_2_nw[8][23]),
    .gather_data_o_8_23                             (gather_data_nw_2_pe[8][23]),
    .gather_valid_o_8_23                            (gather_valid_nw_2_pe[8][23]),
    .gather_ready_i_8_23                            (gather_ready_pe_2_nw[8][23]),
    .cast_data_i_8_24                               (cast_data_pe_2_nw[8][24]),
    .cast_valid_i_8_24                              (cast_valid_pe_2_nw[8][24]),
    .cast_ready_o_8_24                              (cast_ready_nw_2_pe[8][24]),
    .merge_data_i_8_24                              (merge_data_pe_2_nw[8][24]),
    .merge_valid_i_8_24                             (merge_valid_pe_2_nw[8][24]),
    .merge_ready_o_8_24                             (merge_ready_nw_2_pe[8][24]),
    .gather_data_i_8_24                             (gather_data_pe_2_nw[8][24]),
    .gather_valid_i_8_24                            (gather_valid_pe_2_nw[8][24]),
    .gather_ready_o_8_24                            (gather_ready_nw_2_pe[8][24]),

    .cast_data_o_8_24                               (cast_data_nw_2_pe[8][24]),
    .cast_valid_o_8_24                              (cast_valid_nw_2_pe[8][24]),
    .cast_ready_i_8_24                              (cast_ready_pe_2_nw[8][24]),
    .merge_data_o_8_24                              (merge_data_nw_2_pe[8][24]),
    .merge_valid_o_8_24                             (merge_valid_nw_2_pe[8][24]),
    .merge_ready_i_8_24                             (merge_ready_pe_2_nw[8][24]),
    .gather_data_o_8_24                             (gather_data_nw_2_pe[8][24]),
    .gather_valid_o_8_24                            (gather_valid_nw_2_pe[8][24]),
    .gather_ready_i_8_24                            (gather_ready_pe_2_nw[8][24]),
    .cast_data_i_9_0                               (cast_data_pe_2_nw[9][0]),
    .cast_valid_i_9_0                              (cast_valid_pe_2_nw[9][0]),
    .cast_ready_o_9_0                              (cast_ready_nw_2_pe[9][0]),
    .merge_data_i_9_0                              (merge_data_pe_2_nw[9][0]),
    .merge_valid_i_9_0                             (merge_valid_pe_2_nw[9][0]),
    .merge_ready_o_9_0                             (merge_ready_nw_2_pe[9][0]),
    .gather_data_i_9_0                             (gather_data_pe_2_nw[9][0]),
    .gather_valid_i_9_0                            (gather_valid_pe_2_nw[9][0]),
    .gather_ready_o_9_0                            (gather_ready_nw_2_pe[9][0]),

    .cast_data_o_9_0                               (cast_data_nw_2_pe[9][0]),
    .cast_valid_o_9_0                              (cast_valid_nw_2_pe[9][0]),
    .cast_ready_i_9_0                              (cast_ready_pe_2_nw[9][0]),
    .merge_data_o_9_0                              (merge_data_nw_2_pe[9][0]),
    .merge_valid_o_9_0                             (merge_valid_nw_2_pe[9][0]),
    .merge_ready_i_9_0                             (merge_ready_pe_2_nw[9][0]),
    .gather_data_o_9_0                             (gather_data_nw_2_pe[9][0]),
    .gather_valid_o_9_0                            (gather_valid_nw_2_pe[9][0]),
    .gather_ready_i_9_0                            (gather_ready_pe_2_nw[9][0]),
    .cast_data_i_9_1                               (cast_data_pe_2_nw[9][1]),
    .cast_valid_i_9_1                              (cast_valid_pe_2_nw[9][1]),
    .cast_ready_o_9_1                              (cast_ready_nw_2_pe[9][1]),
    .merge_data_i_9_1                              (merge_data_pe_2_nw[9][1]),
    .merge_valid_i_9_1                             (merge_valid_pe_2_nw[9][1]),
    .merge_ready_o_9_1                             (merge_ready_nw_2_pe[9][1]),
    .gather_data_i_9_1                             (gather_data_pe_2_nw[9][1]),
    .gather_valid_i_9_1                            (gather_valid_pe_2_nw[9][1]),
    .gather_ready_o_9_1                            (gather_ready_nw_2_pe[9][1]),

    .cast_data_o_9_1                               (cast_data_nw_2_pe[9][1]),
    .cast_valid_o_9_1                              (cast_valid_nw_2_pe[9][1]),
    .cast_ready_i_9_1                              (cast_ready_pe_2_nw[9][1]),
    .merge_data_o_9_1                              (merge_data_nw_2_pe[9][1]),
    .merge_valid_o_9_1                             (merge_valid_nw_2_pe[9][1]),
    .merge_ready_i_9_1                             (merge_ready_pe_2_nw[9][1]),
    .gather_data_o_9_1                             (gather_data_nw_2_pe[9][1]),
    .gather_valid_o_9_1                            (gather_valid_nw_2_pe[9][1]),
    .gather_ready_i_9_1                            (gather_ready_pe_2_nw[9][1]),
    .cast_data_i_9_2                               (cast_data_pe_2_nw[9][2]),
    .cast_valid_i_9_2                              (cast_valid_pe_2_nw[9][2]),
    .cast_ready_o_9_2                              (cast_ready_nw_2_pe[9][2]),
    .merge_data_i_9_2                              (merge_data_pe_2_nw[9][2]),
    .merge_valid_i_9_2                             (merge_valid_pe_2_nw[9][2]),
    .merge_ready_o_9_2                             (merge_ready_nw_2_pe[9][2]),
    .gather_data_i_9_2                             (gather_data_pe_2_nw[9][2]),
    .gather_valid_i_9_2                            (gather_valid_pe_2_nw[9][2]),
    .gather_ready_o_9_2                            (gather_ready_nw_2_pe[9][2]),

    .cast_data_o_9_2                               (cast_data_nw_2_pe[9][2]),
    .cast_valid_o_9_2                              (cast_valid_nw_2_pe[9][2]),
    .cast_ready_i_9_2                              (cast_ready_pe_2_nw[9][2]),
    .merge_data_o_9_2                              (merge_data_nw_2_pe[9][2]),
    .merge_valid_o_9_2                             (merge_valid_nw_2_pe[9][2]),
    .merge_ready_i_9_2                             (merge_ready_pe_2_nw[9][2]),
    .gather_data_o_9_2                             (gather_data_nw_2_pe[9][2]),
    .gather_valid_o_9_2                            (gather_valid_nw_2_pe[9][2]),
    .gather_ready_i_9_2                            (gather_ready_pe_2_nw[9][2]),
    .cast_data_i_9_3                               (cast_data_pe_2_nw[9][3]),
    .cast_valid_i_9_3                              (cast_valid_pe_2_nw[9][3]),
    .cast_ready_o_9_3                              (cast_ready_nw_2_pe[9][3]),
    .merge_data_i_9_3                              (merge_data_pe_2_nw[9][3]),
    .merge_valid_i_9_3                             (merge_valid_pe_2_nw[9][3]),
    .merge_ready_o_9_3                             (merge_ready_nw_2_pe[9][3]),
    .gather_data_i_9_3                             (gather_data_pe_2_nw[9][3]),
    .gather_valid_i_9_3                            (gather_valid_pe_2_nw[9][3]),
    .gather_ready_o_9_3                            (gather_ready_nw_2_pe[9][3]),

    .cast_data_o_9_3                               (cast_data_nw_2_pe[9][3]),
    .cast_valid_o_9_3                              (cast_valid_nw_2_pe[9][3]),
    .cast_ready_i_9_3                              (cast_ready_pe_2_nw[9][3]),
    .merge_data_o_9_3                              (merge_data_nw_2_pe[9][3]),
    .merge_valid_o_9_3                             (merge_valid_nw_2_pe[9][3]),
    .merge_ready_i_9_3                             (merge_ready_pe_2_nw[9][3]),
    .gather_data_o_9_3                             (gather_data_nw_2_pe[9][3]),
    .gather_valid_o_9_3                            (gather_valid_nw_2_pe[9][3]),
    .gather_ready_i_9_3                            (gather_ready_pe_2_nw[9][3]),
    .cast_data_i_9_4                               (cast_data_pe_2_nw[9][4]),
    .cast_valid_i_9_4                              (cast_valid_pe_2_nw[9][4]),
    .cast_ready_o_9_4                              (cast_ready_nw_2_pe[9][4]),
    .merge_data_i_9_4                              (merge_data_pe_2_nw[9][4]),
    .merge_valid_i_9_4                             (merge_valid_pe_2_nw[9][4]),
    .merge_ready_o_9_4                             (merge_ready_nw_2_pe[9][4]),
    .gather_data_i_9_4                             (gather_data_pe_2_nw[9][4]),
    .gather_valid_i_9_4                            (gather_valid_pe_2_nw[9][4]),
    .gather_ready_o_9_4                            (gather_ready_nw_2_pe[9][4]),

    .cast_data_o_9_4                               (cast_data_nw_2_pe[9][4]),
    .cast_valid_o_9_4                              (cast_valid_nw_2_pe[9][4]),
    .cast_ready_i_9_4                              (cast_ready_pe_2_nw[9][4]),
    .merge_data_o_9_4                              (merge_data_nw_2_pe[9][4]),
    .merge_valid_o_9_4                             (merge_valid_nw_2_pe[9][4]),
    .merge_ready_i_9_4                             (merge_ready_pe_2_nw[9][4]),
    .gather_data_o_9_4                             (gather_data_nw_2_pe[9][4]),
    .gather_valid_o_9_4                            (gather_valid_nw_2_pe[9][4]),
    .gather_ready_i_9_4                            (gather_ready_pe_2_nw[9][4]),
    .cast_data_i_9_5                               (cast_data_pe_2_nw[9][5]),
    .cast_valid_i_9_5                              (cast_valid_pe_2_nw[9][5]),
    .cast_ready_o_9_5                              (cast_ready_nw_2_pe[9][5]),
    .merge_data_i_9_5                              (merge_data_pe_2_nw[9][5]),
    .merge_valid_i_9_5                             (merge_valid_pe_2_nw[9][5]),
    .merge_ready_o_9_5                             (merge_ready_nw_2_pe[9][5]),
    .gather_data_i_9_5                             (gather_data_pe_2_nw[9][5]),
    .gather_valid_i_9_5                            (gather_valid_pe_2_nw[9][5]),
    .gather_ready_o_9_5                            (gather_ready_nw_2_pe[9][5]),

    .cast_data_o_9_5                               (cast_data_nw_2_pe[9][5]),
    .cast_valid_o_9_5                              (cast_valid_nw_2_pe[9][5]),
    .cast_ready_i_9_5                              (cast_ready_pe_2_nw[9][5]),
    .merge_data_o_9_5                              (merge_data_nw_2_pe[9][5]),
    .merge_valid_o_9_5                             (merge_valid_nw_2_pe[9][5]),
    .merge_ready_i_9_5                             (merge_ready_pe_2_nw[9][5]),
    .gather_data_o_9_5                             (gather_data_nw_2_pe[9][5]),
    .gather_valid_o_9_5                            (gather_valid_nw_2_pe[9][5]),
    .gather_ready_i_9_5                            (gather_ready_pe_2_nw[9][5]),
    .cast_data_i_9_6                               (cast_data_pe_2_nw[9][6]),
    .cast_valid_i_9_6                              (cast_valid_pe_2_nw[9][6]),
    .cast_ready_o_9_6                              (cast_ready_nw_2_pe[9][6]),
    .merge_data_i_9_6                              (merge_data_pe_2_nw[9][6]),
    .merge_valid_i_9_6                             (merge_valid_pe_2_nw[9][6]),
    .merge_ready_o_9_6                             (merge_ready_nw_2_pe[9][6]),
    .gather_data_i_9_6                             (gather_data_pe_2_nw[9][6]),
    .gather_valid_i_9_6                            (gather_valid_pe_2_nw[9][6]),
    .gather_ready_o_9_6                            (gather_ready_nw_2_pe[9][6]),

    .cast_data_o_9_6                               (cast_data_nw_2_pe[9][6]),
    .cast_valid_o_9_6                              (cast_valid_nw_2_pe[9][6]),
    .cast_ready_i_9_6                              (cast_ready_pe_2_nw[9][6]),
    .merge_data_o_9_6                              (merge_data_nw_2_pe[9][6]),
    .merge_valid_o_9_6                             (merge_valid_nw_2_pe[9][6]),
    .merge_ready_i_9_6                             (merge_ready_pe_2_nw[9][6]),
    .gather_data_o_9_6                             (gather_data_nw_2_pe[9][6]),
    .gather_valid_o_9_6                            (gather_valid_nw_2_pe[9][6]),
    .gather_ready_i_9_6                            (gather_ready_pe_2_nw[9][6]),
    .cast_data_i_9_7                               (cast_data_pe_2_nw[9][7]),
    .cast_valid_i_9_7                              (cast_valid_pe_2_nw[9][7]),
    .cast_ready_o_9_7                              (cast_ready_nw_2_pe[9][7]),
    .merge_data_i_9_7                              (merge_data_pe_2_nw[9][7]),
    .merge_valid_i_9_7                             (merge_valid_pe_2_nw[9][7]),
    .merge_ready_o_9_7                             (merge_ready_nw_2_pe[9][7]),
    .gather_data_i_9_7                             (gather_data_pe_2_nw[9][7]),
    .gather_valid_i_9_7                            (gather_valid_pe_2_nw[9][7]),
    .gather_ready_o_9_7                            (gather_ready_nw_2_pe[9][7]),

    .cast_data_o_9_7                               (cast_data_nw_2_pe[9][7]),
    .cast_valid_o_9_7                              (cast_valid_nw_2_pe[9][7]),
    .cast_ready_i_9_7                              (cast_ready_pe_2_nw[9][7]),
    .merge_data_o_9_7                              (merge_data_nw_2_pe[9][7]),
    .merge_valid_o_9_7                             (merge_valid_nw_2_pe[9][7]),
    .merge_ready_i_9_7                             (merge_ready_pe_2_nw[9][7]),
    .gather_data_o_9_7                             (gather_data_nw_2_pe[9][7]),
    .gather_valid_o_9_7                            (gather_valid_nw_2_pe[9][7]),
    .gather_ready_i_9_7                            (gather_ready_pe_2_nw[9][7]),
    .cast_data_i_9_8                               (cast_data_pe_2_nw[9][8]),
    .cast_valid_i_9_8                              (cast_valid_pe_2_nw[9][8]),
    .cast_ready_o_9_8                              (cast_ready_nw_2_pe[9][8]),
    .merge_data_i_9_8                              (merge_data_pe_2_nw[9][8]),
    .merge_valid_i_9_8                             (merge_valid_pe_2_nw[9][8]),
    .merge_ready_o_9_8                             (merge_ready_nw_2_pe[9][8]),
    .gather_data_i_9_8                             (gather_data_pe_2_nw[9][8]),
    .gather_valid_i_9_8                            (gather_valid_pe_2_nw[9][8]),
    .gather_ready_o_9_8                            (gather_ready_nw_2_pe[9][8]),

    .cast_data_o_9_8                               (cast_data_nw_2_pe[9][8]),
    .cast_valid_o_9_8                              (cast_valid_nw_2_pe[9][8]),
    .cast_ready_i_9_8                              (cast_ready_pe_2_nw[9][8]),
    .merge_data_o_9_8                              (merge_data_nw_2_pe[9][8]),
    .merge_valid_o_9_8                             (merge_valid_nw_2_pe[9][8]),
    .merge_ready_i_9_8                             (merge_ready_pe_2_nw[9][8]),
    .gather_data_o_9_8                             (gather_data_nw_2_pe[9][8]),
    .gather_valid_o_9_8                            (gather_valid_nw_2_pe[9][8]),
    .gather_ready_i_9_8                            (gather_ready_pe_2_nw[9][8]),
    .cast_data_i_9_9                               (cast_data_pe_2_nw[9][9]),
    .cast_valid_i_9_9                              (cast_valid_pe_2_nw[9][9]),
    .cast_ready_o_9_9                              (cast_ready_nw_2_pe[9][9]),
    .merge_data_i_9_9                              (merge_data_pe_2_nw[9][9]),
    .merge_valid_i_9_9                             (merge_valid_pe_2_nw[9][9]),
    .merge_ready_o_9_9                             (merge_ready_nw_2_pe[9][9]),
    .gather_data_i_9_9                             (gather_data_pe_2_nw[9][9]),
    .gather_valid_i_9_9                            (gather_valid_pe_2_nw[9][9]),
    .gather_ready_o_9_9                            (gather_ready_nw_2_pe[9][9]),

    .cast_data_o_9_9                               (cast_data_nw_2_pe[9][9]),
    .cast_valid_o_9_9                              (cast_valid_nw_2_pe[9][9]),
    .cast_ready_i_9_9                              (cast_ready_pe_2_nw[9][9]),
    .merge_data_o_9_9                              (merge_data_nw_2_pe[9][9]),
    .merge_valid_o_9_9                             (merge_valid_nw_2_pe[9][9]),
    .merge_ready_i_9_9                             (merge_ready_pe_2_nw[9][9]),
    .gather_data_o_9_9                             (gather_data_nw_2_pe[9][9]),
    .gather_valid_o_9_9                            (gather_valid_nw_2_pe[9][9]),
    .gather_ready_i_9_9                            (gather_ready_pe_2_nw[9][9]),
    .cast_data_i_9_10                               (cast_data_pe_2_nw[9][10]),
    .cast_valid_i_9_10                              (cast_valid_pe_2_nw[9][10]),
    .cast_ready_o_9_10                              (cast_ready_nw_2_pe[9][10]),
    .merge_data_i_9_10                              (merge_data_pe_2_nw[9][10]),
    .merge_valid_i_9_10                             (merge_valid_pe_2_nw[9][10]),
    .merge_ready_o_9_10                             (merge_ready_nw_2_pe[9][10]),
    .gather_data_i_9_10                             (gather_data_pe_2_nw[9][10]),
    .gather_valid_i_9_10                            (gather_valid_pe_2_nw[9][10]),
    .gather_ready_o_9_10                            (gather_ready_nw_2_pe[9][10]),

    .cast_data_o_9_10                               (cast_data_nw_2_pe[9][10]),
    .cast_valid_o_9_10                              (cast_valid_nw_2_pe[9][10]),
    .cast_ready_i_9_10                              (cast_ready_pe_2_nw[9][10]),
    .merge_data_o_9_10                              (merge_data_nw_2_pe[9][10]),
    .merge_valid_o_9_10                             (merge_valid_nw_2_pe[9][10]),
    .merge_ready_i_9_10                             (merge_ready_pe_2_nw[9][10]),
    .gather_data_o_9_10                             (gather_data_nw_2_pe[9][10]),
    .gather_valid_o_9_10                            (gather_valid_nw_2_pe[9][10]),
    .gather_ready_i_9_10                            (gather_ready_pe_2_nw[9][10]),
    .cast_data_i_9_11                               (cast_data_pe_2_nw[9][11]),
    .cast_valid_i_9_11                              (cast_valid_pe_2_nw[9][11]),
    .cast_ready_o_9_11                              (cast_ready_nw_2_pe[9][11]),
    .merge_data_i_9_11                              (merge_data_pe_2_nw[9][11]),
    .merge_valid_i_9_11                             (merge_valid_pe_2_nw[9][11]),
    .merge_ready_o_9_11                             (merge_ready_nw_2_pe[9][11]),
    .gather_data_i_9_11                             (gather_data_pe_2_nw[9][11]),
    .gather_valid_i_9_11                            (gather_valid_pe_2_nw[9][11]),
    .gather_ready_o_9_11                            (gather_ready_nw_2_pe[9][11]),

    .cast_data_o_9_11                               (cast_data_nw_2_pe[9][11]),
    .cast_valid_o_9_11                              (cast_valid_nw_2_pe[9][11]),
    .cast_ready_i_9_11                              (cast_ready_pe_2_nw[9][11]),
    .merge_data_o_9_11                              (merge_data_nw_2_pe[9][11]),
    .merge_valid_o_9_11                             (merge_valid_nw_2_pe[9][11]),
    .merge_ready_i_9_11                             (merge_ready_pe_2_nw[9][11]),
    .gather_data_o_9_11                             (gather_data_nw_2_pe[9][11]),
    .gather_valid_o_9_11                            (gather_valid_nw_2_pe[9][11]),
    .gather_ready_i_9_11                            (gather_ready_pe_2_nw[9][11]),
    .cast_data_i_9_12                               (cast_data_pe_2_nw[9][12]),
    .cast_valid_i_9_12                              (cast_valid_pe_2_nw[9][12]),
    .cast_ready_o_9_12                              (cast_ready_nw_2_pe[9][12]),
    .merge_data_i_9_12                              (merge_data_pe_2_nw[9][12]),
    .merge_valid_i_9_12                             (merge_valid_pe_2_nw[9][12]),
    .merge_ready_o_9_12                             (merge_ready_nw_2_pe[9][12]),
    .gather_data_i_9_12                             (gather_data_pe_2_nw[9][12]),
    .gather_valid_i_9_12                            (gather_valid_pe_2_nw[9][12]),
    .gather_ready_o_9_12                            (gather_ready_nw_2_pe[9][12]),

    .cast_data_o_9_12                               (cast_data_nw_2_pe[9][12]),
    .cast_valid_o_9_12                              (cast_valid_nw_2_pe[9][12]),
    .cast_ready_i_9_12                              (cast_ready_pe_2_nw[9][12]),
    .merge_data_o_9_12                              (merge_data_nw_2_pe[9][12]),
    .merge_valid_o_9_12                             (merge_valid_nw_2_pe[9][12]),
    .merge_ready_i_9_12                             (merge_ready_pe_2_nw[9][12]),
    .gather_data_o_9_12                             (gather_data_nw_2_pe[9][12]),
    .gather_valid_o_9_12                            (gather_valid_nw_2_pe[9][12]),
    .gather_ready_i_9_12                            (gather_ready_pe_2_nw[9][12]),
    .cast_data_i_9_13                               (cast_data_pe_2_nw[9][13]),
    .cast_valid_i_9_13                              (cast_valid_pe_2_nw[9][13]),
    .cast_ready_o_9_13                              (cast_ready_nw_2_pe[9][13]),
    .merge_data_i_9_13                              (merge_data_pe_2_nw[9][13]),
    .merge_valid_i_9_13                             (merge_valid_pe_2_nw[9][13]),
    .merge_ready_o_9_13                             (merge_ready_nw_2_pe[9][13]),
    .gather_data_i_9_13                             (gather_data_pe_2_nw[9][13]),
    .gather_valid_i_9_13                            (gather_valid_pe_2_nw[9][13]),
    .gather_ready_o_9_13                            (gather_ready_nw_2_pe[9][13]),

    .cast_data_o_9_13                               (cast_data_nw_2_pe[9][13]),
    .cast_valid_o_9_13                              (cast_valid_nw_2_pe[9][13]),
    .cast_ready_i_9_13                              (cast_ready_pe_2_nw[9][13]),
    .merge_data_o_9_13                              (merge_data_nw_2_pe[9][13]),
    .merge_valid_o_9_13                             (merge_valid_nw_2_pe[9][13]),
    .merge_ready_i_9_13                             (merge_ready_pe_2_nw[9][13]),
    .gather_data_o_9_13                             (gather_data_nw_2_pe[9][13]),
    .gather_valid_o_9_13                            (gather_valid_nw_2_pe[9][13]),
    .gather_ready_i_9_13                            (gather_ready_pe_2_nw[9][13]),
    .cast_data_i_9_14                               (cast_data_pe_2_nw[9][14]),
    .cast_valid_i_9_14                              (cast_valid_pe_2_nw[9][14]),
    .cast_ready_o_9_14                              (cast_ready_nw_2_pe[9][14]),
    .merge_data_i_9_14                              (merge_data_pe_2_nw[9][14]),
    .merge_valid_i_9_14                             (merge_valid_pe_2_nw[9][14]),
    .merge_ready_o_9_14                             (merge_ready_nw_2_pe[9][14]),
    .gather_data_i_9_14                             (gather_data_pe_2_nw[9][14]),
    .gather_valid_i_9_14                            (gather_valid_pe_2_nw[9][14]),
    .gather_ready_o_9_14                            (gather_ready_nw_2_pe[9][14]),

    .cast_data_o_9_14                               (cast_data_nw_2_pe[9][14]),
    .cast_valid_o_9_14                              (cast_valid_nw_2_pe[9][14]),
    .cast_ready_i_9_14                              (cast_ready_pe_2_nw[9][14]),
    .merge_data_o_9_14                              (merge_data_nw_2_pe[9][14]),
    .merge_valid_o_9_14                             (merge_valid_nw_2_pe[9][14]),
    .merge_ready_i_9_14                             (merge_ready_pe_2_nw[9][14]),
    .gather_data_o_9_14                             (gather_data_nw_2_pe[9][14]),
    .gather_valid_o_9_14                            (gather_valid_nw_2_pe[9][14]),
    .gather_ready_i_9_14                            (gather_ready_pe_2_nw[9][14]),
    .cast_data_i_9_15                               (cast_data_pe_2_nw[9][15]),
    .cast_valid_i_9_15                              (cast_valid_pe_2_nw[9][15]),
    .cast_ready_o_9_15                              (cast_ready_nw_2_pe[9][15]),
    .merge_data_i_9_15                              (merge_data_pe_2_nw[9][15]),
    .merge_valid_i_9_15                             (merge_valid_pe_2_nw[9][15]),
    .merge_ready_o_9_15                             (merge_ready_nw_2_pe[9][15]),
    .gather_data_i_9_15                             (gather_data_pe_2_nw[9][15]),
    .gather_valid_i_9_15                            (gather_valid_pe_2_nw[9][15]),
    .gather_ready_o_9_15                            (gather_ready_nw_2_pe[9][15]),

    .cast_data_o_9_15                               (cast_data_nw_2_pe[9][15]),
    .cast_valid_o_9_15                              (cast_valid_nw_2_pe[9][15]),
    .cast_ready_i_9_15                              (cast_ready_pe_2_nw[9][15]),
    .merge_data_o_9_15                              (merge_data_nw_2_pe[9][15]),
    .merge_valid_o_9_15                             (merge_valid_nw_2_pe[9][15]),
    .merge_ready_i_9_15                             (merge_ready_pe_2_nw[9][15]),
    .gather_data_o_9_15                             (gather_data_nw_2_pe[9][15]),
    .gather_valid_o_9_15                            (gather_valid_nw_2_pe[9][15]),
    .gather_ready_i_9_15                            (gather_ready_pe_2_nw[9][15]),
    .cast_data_i_9_16                               (cast_data_pe_2_nw[9][16]),
    .cast_valid_i_9_16                              (cast_valid_pe_2_nw[9][16]),
    .cast_ready_o_9_16                              (cast_ready_nw_2_pe[9][16]),
    .merge_data_i_9_16                              (merge_data_pe_2_nw[9][16]),
    .merge_valid_i_9_16                             (merge_valid_pe_2_nw[9][16]),
    .merge_ready_o_9_16                             (merge_ready_nw_2_pe[9][16]),
    .gather_data_i_9_16                             (gather_data_pe_2_nw[9][16]),
    .gather_valid_i_9_16                            (gather_valid_pe_2_nw[9][16]),
    .gather_ready_o_9_16                            (gather_ready_nw_2_pe[9][16]),

    .cast_data_o_9_16                               (cast_data_nw_2_pe[9][16]),
    .cast_valid_o_9_16                              (cast_valid_nw_2_pe[9][16]),
    .cast_ready_i_9_16                              (cast_ready_pe_2_nw[9][16]),
    .merge_data_o_9_16                              (merge_data_nw_2_pe[9][16]),
    .merge_valid_o_9_16                             (merge_valid_nw_2_pe[9][16]),
    .merge_ready_i_9_16                             (merge_ready_pe_2_nw[9][16]),
    .gather_data_o_9_16                             (gather_data_nw_2_pe[9][16]),
    .gather_valid_o_9_16                            (gather_valid_nw_2_pe[9][16]),
    .gather_ready_i_9_16                            (gather_ready_pe_2_nw[9][16]),
    .cast_data_i_9_17                               (cast_data_pe_2_nw[9][17]),
    .cast_valid_i_9_17                              (cast_valid_pe_2_nw[9][17]),
    .cast_ready_o_9_17                              (cast_ready_nw_2_pe[9][17]),
    .merge_data_i_9_17                              (merge_data_pe_2_nw[9][17]),
    .merge_valid_i_9_17                             (merge_valid_pe_2_nw[9][17]),
    .merge_ready_o_9_17                             (merge_ready_nw_2_pe[9][17]),
    .gather_data_i_9_17                             (gather_data_pe_2_nw[9][17]),
    .gather_valid_i_9_17                            (gather_valid_pe_2_nw[9][17]),
    .gather_ready_o_9_17                            (gather_ready_nw_2_pe[9][17]),

    .cast_data_o_9_17                               (cast_data_nw_2_pe[9][17]),
    .cast_valid_o_9_17                              (cast_valid_nw_2_pe[9][17]),
    .cast_ready_i_9_17                              (cast_ready_pe_2_nw[9][17]),
    .merge_data_o_9_17                              (merge_data_nw_2_pe[9][17]),
    .merge_valid_o_9_17                             (merge_valid_nw_2_pe[9][17]),
    .merge_ready_i_9_17                             (merge_ready_pe_2_nw[9][17]),
    .gather_data_o_9_17                             (gather_data_nw_2_pe[9][17]),
    .gather_valid_o_9_17                            (gather_valid_nw_2_pe[9][17]),
    .gather_ready_i_9_17                            (gather_ready_pe_2_nw[9][17]),
    .cast_data_i_9_18                               (cast_data_pe_2_nw[9][18]),
    .cast_valid_i_9_18                              (cast_valid_pe_2_nw[9][18]),
    .cast_ready_o_9_18                              (cast_ready_nw_2_pe[9][18]),
    .merge_data_i_9_18                              (merge_data_pe_2_nw[9][18]),
    .merge_valid_i_9_18                             (merge_valid_pe_2_nw[9][18]),
    .merge_ready_o_9_18                             (merge_ready_nw_2_pe[9][18]),
    .gather_data_i_9_18                             (gather_data_pe_2_nw[9][18]),
    .gather_valid_i_9_18                            (gather_valid_pe_2_nw[9][18]),
    .gather_ready_o_9_18                            (gather_ready_nw_2_pe[9][18]),

    .cast_data_o_9_18                               (cast_data_nw_2_pe[9][18]),
    .cast_valid_o_9_18                              (cast_valid_nw_2_pe[9][18]),
    .cast_ready_i_9_18                              (cast_ready_pe_2_nw[9][18]),
    .merge_data_o_9_18                              (merge_data_nw_2_pe[9][18]),
    .merge_valid_o_9_18                             (merge_valid_nw_2_pe[9][18]),
    .merge_ready_i_9_18                             (merge_ready_pe_2_nw[9][18]),
    .gather_data_o_9_18                             (gather_data_nw_2_pe[9][18]),
    .gather_valid_o_9_18                            (gather_valid_nw_2_pe[9][18]),
    .gather_ready_i_9_18                            (gather_ready_pe_2_nw[9][18]),
    .cast_data_i_9_19                               (cast_data_pe_2_nw[9][19]),
    .cast_valid_i_9_19                              (cast_valid_pe_2_nw[9][19]),
    .cast_ready_o_9_19                              (cast_ready_nw_2_pe[9][19]),
    .merge_data_i_9_19                              (merge_data_pe_2_nw[9][19]),
    .merge_valid_i_9_19                             (merge_valid_pe_2_nw[9][19]),
    .merge_ready_o_9_19                             (merge_ready_nw_2_pe[9][19]),
    .gather_data_i_9_19                             (gather_data_pe_2_nw[9][19]),
    .gather_valid_i_9_19                            (gather_valid_pe_2_nw[9][19]),
    .gather_ready_o_9_19                            (gather_ready_nw_2_pe[9][19]),

    .cast_data_o_9_19                               (cast_data_nw_2_pe[9][19]),
    .cast_valid_o_9_19                              (cast_valid_nw_2_pe[9][19]),
    .cast_ready_i_9_19                              (cast_ready_pe_2_nw[9][19]),
    .merge_data_o_9_19                              (merge_data_nw_2_pe[9][19]),
    .merge_valid_o_9_19                             (merge_valid_nw_2_pe[9][19]),
    .merge_ready_i_9_19                             (merge_ready_pe_2_nw[9][19]),
    .gather_data_o_9_19                             (gather_data_nw_2_pe[9][19]),
    .gather_valid_o_9_19                            (gather_valid_nw_2_pe[9][19]),
    .gather_ready_i_9_19                            (gather_ready_pe_2_nw[9][19]),
    .cast_data_i_9_20                               (cast_data_pe_2_nw[9][20]),
    .cast_valid_i_9_20                              (cast_valid_pe_2_nw[9][20]),
    .cast_ready_o_9_20                              (cast_ready_nw_2_pe[9][20]),
    .merge_data_i_9_20                              (merge_data_pe_2_nw[9][20]),
    .merge_valid_i_9_20                             (merge_valid_pe_2_nw[9][20]),
    .merge_ready_o_9_20                             (merge_ready_nw_2_pe[9][20]),
    .gather_data_i_9_20                             (gather_data_pe_2_nw[9][20]),
    .gather_valid_i_9_20                            (gather_valid_pe_2_nw[9][20]),
    .gather_ready_o_9_20                            (gather_ready_nw_2_pe[9][20]),

    .cast_data_o_9_20                               (cast_data_nw_2_pe[9][20]),
    .cast_valid_o_9_20                              (cast_valid_nw_2_pe[9][20]),
    .cast_ready_i_9_20                              (cast_ready_pe_2_nw[9][20]),
    .merge_data_o_9_20                              (merge_data_nw_2_pe[9][20]),
    .merge_valid_o_9_20                             (merge_valid_nw_2_pe[9][20]),
    .merge_ready_i_9_20                             (merge_ready_pe_2_nw[9][20]),
    .gather_data_o_9_20                             (gather_data_nw_2_pe[9][20]),
    .gather_valid_o_9_20                            (gather_valid_nw_2_pe[9][20]),
    .gather_ready_i_9_20                            (gather_ready_pe_2_nw[9][20]),
    .cast_data_i_9_21                               (cast_data_pe_2_nw[9][21]),
    .cast_valid_i_9_21                              (cast_valid_pe_2_nw[9][21]),
    .cast_ready_o_9_21                              (cast_ready_nw_2_pe[9][21]),
    .merge_data_i_9_21                              (merge_data_pe_2_nw[9][21]),
    .merge_valid_i_9_21                             (merge_valid_pe_2_nw[9][21]),
    .merge_ready_o_9_21                             (merge_ready_nw_2_pe[9][21]),
    .gather_data_i_9_21                             (gather_data_pe_2_nw[9][21]),
    .gather_valid_i_9_21                            (gather_valid_pe_2_nw[9][21]),
    .gather_ready_o_9_21                            (gather_ready_nw_2_pe[9][21]),

    .cast_data_o_9_21                               (cast_data_nw_2_pe[9][21]),
    .cast_valid_o_9_21                              (cast_valid_nw_2_pe[9][21]),
    .cast_ready_i_9_21                              (cast_ready_pe_2_nw[9][21]),
    .merge_data_o_9_21                              (merge_data_nw_2_pe[9][21]),
    .merge_valid_o_9_21                             (merge_valid_nw_2_pe[9][21]),
    .merge_ready_i_9_21                             (merge_ready_pe_2_nw[9][21]),
    .gather_data_o_9_21                             (gather_data_nw_2_pe[9][21]),
    .gather_valid_o_9_21                            (gather_valid_nw_2_pe[9][21]),
    .gather_ready_i_9_21                            (gather_ready_pe_2_nw[9][21]),
    .cast_data_i_9_22                               (cast_data_pe_2_nw[9][22]),
    .cast_valid_i_9_22                              (cast_valid_pe_2_nw[9][22]),
    .cast_ready_o_9_22                              (cast_ready_nw_2_pe[9][22]),
    .merge_data_i_9_22                              (merge_data_pe_2_nw[9][22]),
    .merge_valid_i_9_22                             (merge_valid_pe_2_nw[9][22]),
    .merge_ready_o_9_22                             (merge_ready_nw_2_pe[9][22]),
    .gather_data_i_9_22                             (gather_data_pe_2_nw[9][22]),
    .gather_valid_i_9_22                            (gather_valid_pe_2_nw[9][22]),
    .gather_ready_o_9_22                            (gather_ready_nw_2_pe[9][22]),

    .cast_data_o_9_22                               (cast_data_nw_2_pe[9][22]),
    .cast_valid_o_9_22                              (cast_valid_nw_2_pe[9][22]),
    .cast_ready_i_9_22                              (cast_ready_pe_2_nw[9][22]),
    .merge_data_o_9_22                              (merge_data_nw_2_pe[9][22]),
    .merge_valid_o_9_22                             (merge_valid_nw_2_pe[9][22]),
    .merge_ready_i_9_22                             (merge_ready_pe_2_nw[9][22]),
    .gather_data_o_9_22                             (gather_data_nw_2_pe[9][22]),
    .gather_valid_o_9_22                            (gather_valid_nw_2_pe[9][22]),
    .gather_ready_i_9_22                            (gather_ready_pe_2_nw[9][22]),
    .cast_data_i_9_23                               (cast_data_pe_2_nw[9][23]),
    .cast_valid_i_9_23                              (cast_valid_pe_2_nw[9][23]),
    .cast_ready_o_9_23                              (cast_ready_nw_2_pe[9][23]),
    .merge_data_i_9_23                              (merge_data_pe_2_nw[9][23]),
    .merge_valid_i_9_23                             (merge_valid_pe_2_nw[9][23]),
    .merge_ready_o_9_23                             (merge_ready_nw_2_pe[9][23]),
    .gather_data_i_9_23                             (gather_data_pe_2_nw[9][23]),
    .gather_valid_i_9_23                            (gather_valid_pe_2_nw[9][23]),
    .gather_ready_o_9_23                            (gather_ready_nw_2_pe[9][23]),

    .cast_data_o_9_23                               (cast_data_nw_2_pe[9][23]),
    .cast_valid_o_9_23                              (cast_valid_nw_2_pe[9][23]),
    .cast_ready_i_9_23                              (cast_ready_pe_2_nw[9][23]),
    .merge_data_o_9_23                              (merge_data_nw_2_pe[9][23]),
    .merge_valid_o_9_23                             (merge_valid_nw_2_pe[9][23]),
    .merge_ready_i_9_23                             (merge_ready_pe_2_nw[9][23]),
    .gather_data_o_9_23                             (gather_data_nw_2_pe[9][23]),
    .gather_valid_o_9_23                            (gather_valid_nw_2_pe[9][23]),
    .gather_ready_i_9_23                            (gather_ready_pe_2_nw[9][23]),
    .cast_data_i_9_24                               (cast_data_pe_2_nw[9][24]),
    .cast_valid_i_9_24                              (cast_valid_pe_2_nw[9][24]),
    .cast_ready_o_9_24                              (cast_ready_nw_2_pe[9][24]),
    .merge_data_i_9_24                              (merge_data_pe_2_nw[9][24]),
    .merge_valid_i_9_24                             (merge_valid_pe_2_nw[9][24]),
    .merge_ready_o_9_24                             (merge_ready_nw_2_pe[9][24]),
    .gather_data_i_9_24                             (gather_data_pe_2_nw[9][24]),
    .gather_valid_i_9_24                            (gather_valid_pe_2_nw[9][24]),
    .gather_ready_o_9_24                            (gather_ready_nw_2_pe[9][24]),

    .cast_data_o_9_24                               (cast_data_nw_2_pe[9][24]),
    .cast_valid_o_9_24                              (cast_valid_nw_2_pe[9][24]),
    .cast_ready_i_9_24                              (cast_ready_pe_2_nw[9][24]),
    .merge_data_o_9_24                              (merge_data_nw_2_pe[9][24]),
    .merge_valid_o_9_24                             (merge_valid_nw_2_pe[9][24]),
    .merge_ready_i_9_24                             (merge_ready_pe_2_nw[9][24]),
    .gather_data_o_9_24                             (gather_data_nw_2_pe[9][24]),
    .gather_valid_o_9_24                            (gather_valid_nw_2_pe[9][24]),
    .gather_ready_i_9_24                            (gather_ready_pe_2_nw[9][24])
);

virtual_pe #(
    .cast_out                                          (cast_out_0_0),
    .merge_in                                          (merge_in_0_0),
    .merge_out                                         (merge_out_0_0),
    .gather_in                                         (gather_in_0_0),
    .gather_out                                        (gather_out_0_0),
    .x                                                 (0),
    .y                                                 (0)
)vpe_0_0(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[0][0]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[0][0]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[0][0]),
    .cast_data_o                                       (cast_data_pe_2_nw[0][0]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[0][0]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[0][0]),
    .merge_data_i                                      (merge_data_nw_2_pe[0][0]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[0][0]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[0][0]),
    .merge_data_o                                      (merge_data_pe_2_nw[0][0]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[0][0]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[0][0]),
    .gather_data_i                                     (gather_data_nw_2_pe[0][0]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[0][0]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[0][0]),
    .gather_data_o                                     (gather_data_pe_2_nw[0][0]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[0][0]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[0][0])
);


virtual_pe #(
    .cast_out                                          (cast_out_0_1),
    .merge_in                                          (merge_in_0_1),
    .merge_out                                         (merge_out_0_1),
    .gather_in                                         (gather_in_0_1),
    .gather_out                                        (gather_out_0_1),
    .x                                                 (0),
    .y                                                 (1)
)vpe_0_1(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[0][1]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[0][1]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[0][1]),
    .cast_data_o                                       (cast_data_pe_2_nw[0][1]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[0][1]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[0][1]),
    .merge_data_i                                      (merge_data_nw_2_pe[0][1]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[0][1]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[0][1]),
    .merge_data_o                                      (merge_data_pe_2_nw[0][1]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[0][1]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[0][1]),
    .gather_data_i                                     (gather_data_nw_2_pe[0][1]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[0][1]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[0][1]),
    .gather_data_o                                     (gather_data_pe_2_nw[0][1]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[0][1]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[0][1])
);


virtual_pe #(
    .cast_out                                          (cast_out_0_2),
    .merge_in                                          (merge_in_0_2),
    .merge_out                                         (merge_out_0_2),
    .gather_in                                         (gather_in_0_2),
    .gather_out                                        (gather_out_0_2),
    .x                                                 (0),
    .y                                                 (2)
)vpe_0_2(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[0][2]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[0][2]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[0][2]),
    .cast_data_o                                       (cast_data_pe_2_nw[0][2]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[0][2]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[0][2]),
    .merge_data_i                                      (merge_data_nw_2_pe[0][2]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[0][2]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[0][2]),
    .merge_data_o                                      (merge_data_pe_2_nw[0][2]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[0][2]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[0][2]),
    .gather_data_i                                     (gather_data_nw_2_pe[0][2]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[0][2]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[0][2]),
    .gather_data_o                                     (gather_data_pe_2_nw[0][2]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[0][2]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[0][2])
);


virtual_pe #(
    .cast_out                                          (cast_out_0_3),
    .merge_in                                          (merge_in_0_3),
    .merge_out                                         (merge_out_0_3),
    .gather_in                                         (gather_in_0_3),
    .gather_out                                        (gather_out_0_3),
    .x                                                 (0),
    .y                                                 (3)
)vpe_0_3(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[0][3]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[0][3]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[0][3]),
    .cast_data_o                                       (cast_data_pe_2_nw[0][3]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[0][3]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[0][3]),
    .merge_data_i                                      (merge_data_nw_2_pe[0][3]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[0][3]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[0][3]),
    .merge_data_o                                      (merge_data_pe_2_nw[0][3]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[0][3]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[0][3]),
    .gather_data_i                                     (gather_data_nw_2_pe[0][3]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[0][3]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[0][3]),
    .gather_data_o                                     (gather_data_pe_2_nw[0][3]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[0][3]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[0][3])
);


virtual_pe #(
    .cast_out                                          (cast_out_0_4),
    .merge_in                                          (merge_in_0_4),
    .merge_out                                         (merge_out_0_4),
    .gather_in                                         (gather_in_0_4),
    .gather_out                                        (gather_out_0_4),
    .x                                                 (0),
    .y                                                 (4)
)vpe_0_4(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[0][4]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[0][4]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[0][4]),
    .cast_data_o                                       (cast_data_pe_2_nw[0][4]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[0][4]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[0][4]),
    .merge_data_i                                      (merge_data_nw_2_pe[0][4]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[0][4]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[0][4]),
    .merge_data_o                                      (merge_data_pe_2_nw[0][4]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[0][4]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[0][4]),
    .gather_data_i                                     (gather_data_nw_2_pe[0][4]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[0][4]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[0][4]),
    .gather_data_o                                     (gather_data_pe_2_nw[0][4]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[0][4]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[0][4])
);


virtual_pe #(
    .cast_out                                          (cast_out_0_5),
    .merge_in                                          (merge_in_0_5),
    .merge_out                                         (merge_out_0_5),
    .gather_in                                         (gather_in_0_5),
    .gather_out                                        (gather_out_0_5),
    .x                                                 (0),
    .y                                                 (5)
)vpe_0_5(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[0][5]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[0][5]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[0][5]),
    .cast_data_o                                       (cast_data_pe_2_nw[0][5]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[0][5]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[0][5]),
    .merge_data_i                                      (merge_data_nw_2_pe[0][5]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[0][5]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[0][5]),
    .merge_data_o                                      (merge_data_pe_2_nw[0][5]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[0][5]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[0][5]),
    .gather_data_i                                     (gather_data_nw_2_pe[0][5]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[0][5]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[0][5]),
    .gather_data_o                                     (gather_data_pe_2_nw[0][5]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[0][5]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[0][5])
);


virtual_pe #(
    .cast_out                                          (cast_out_0_6),
    .merge_in                                          (merge_in_0_6),
    .merge_out                                         (merge_out_0_6),
    .gather_in                                         (gather_in_0_6),
    .gather_out                                        (gather_out_0_6),
    .x                                                 (0),
    .y                                                 (6)
)vpe_0_6(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[0][6]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[0][6]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[0][6]),
    .cast_data_o                                       (cast_data_pe_2_nw[0][6]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[0][6]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[0][6]),
    .merge_data_i                                      (merge_data_nw_2_pe[0][6]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[0][6]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[0][6]),
    .merge_data_o                                      (merge_data_pe_2_nw[0][6]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[0][6]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[0][6]),
    .gather_data_i                                     (gather_data_nw_2_pe[0][6]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[0][6]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[0][6]),
    .gather_data_o                                     (gather_data_pe_2_nw[0][6]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[0][6]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[0][6])
);


virtual_pe #(
    .cast_out                                          (cast_out_0_7),
    .merge_in                                          (merge_in_0_7),
    .merge_out                                         (merge_out_0_7),
    .gather_in                                         (gather_in_0_7),
    .gather_out                                        (gather_out_0_7),
    .x                                                 (0),
    .y                                                 (7)
)vpe_0_7(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[0][7]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[0][7]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[0][7]),
    .cast_data_o                                       (cast_data_pe_2_nw[0][7]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[0][7]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[0][7]),
    .merge_data_i                                      (merge_data_nw_2_pe[0][7]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[0][7]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[0][7]),
    .merge_data_o                                      (merge_data_pe_2_nw[0][7]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[0][7]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[0][7]),
    .gather_data_i                                     (gather_data_nw_2_pe[0][7]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[0][7]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[0][7]),
    .gather_data_o                                     (gather_data_pe_2_nw[0][7]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[0][7]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[0][7])
);


virtual_pe #(
    .cast_out                                          (cast_out_0_8),
    .merge_in                                          (merge_in_0_8),
    .merge_out                                         (merge_out_0_8),
    .gather_in                                         (gather_in_0_8),
    .gather_out                                        (gather_out_0_8),
    .x                                                 (0),
    .y                                                 (8)
)vpe_0_8(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[0][8]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[0][8]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[0][8]),
    .cast_data_o                                       (cast_data_pe_2_nw[0][8]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[0][8]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[0][8]),
    .merge_data_i                                      (merge_data_nw_2_pe[0][8]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[0][8]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[0][8]),
    .merge_data_o                                      (merge_data_pe_2_nw[0][8]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[0][8]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[0][8]),
    .gather_data_i                                     (gather_data_nw_2_pe[0][8]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[0][8]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[0][8]),
    .gather_data_o                                     (gather_data_pe_2_nw[0][8]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[0][8]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[0][8])
);


virtual_pe #(
    .cast_out                                          (cast_out_0_9),
    .merge_in                                          (merge_in_0_9),
    .merge_out                                         (merge_out_0_9),
    .gather_in                                         (gather_in_0_9),
    .gather_out                                        (gather_out_0_9),
    .x                                                 (0),
    .y                                                 (9)
)vpe_0_9(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[0][9]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[0][9]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[0][9]),
    .cast_data_o                                       (cast_data_pe_2_nw[0][9]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[0][9]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[0][9]),
    .merge_data_i                                      (merge_data_nw_2_pe[0][9]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[0][9]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[0][9]),
    .merge_data_o                                      (merge_data_pe_2_nw[0][9]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[0][9]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[0][9]),
    .gather_data_i                                     (gather_data_nw_2_pe[0][9]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[0][9]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[0][9]),
    .gather_data_o                                     (gather_data_pe_2_nw[0][9]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[0][9]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[0][9])
);


virtual_pe #(
    .cast_out                                          (cast_out_0_10),
    .merge_in                                          (merge_in_0_10),
    .merge_out                                         (merge_out_0_10),
    .gather_in                                         (gather_in_0_10),
    .gather_out                                        (gather_out_0_10),
    .x                                                 (0),
    .y                                                 (10)
)vpe_0_10(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[0][10]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[0][10]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[0][10]),
    .cast_data_o                                       (cast_data_pe_2_nw[0][10]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[0][10]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[0][10]),
    .merge_data_i                                      (merge_data_nw_2_pe[0][10]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[0][10]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[0][10]),
    .merge_data_o                                      (merge_data_pe_2_nw[0][10]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[0][10]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[0][10]),
    .gather_data_i                                     (gather_data_nw_2_pe[0][10]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[0][10]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[0][10]),
    .gather_data_o                                     (gather_data_pe_2_nw[0][10]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[0][10]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[0][10])
);


virtual_pe #(
    .cast_out                                          (cast_out_0_11),
    .merge_in                                          (merge_in_0_11),
    .merge_out                                         (merge_out_0_11),
    .gather_in                                         (gather_in_0_11),
    .gather_out                                        (gather_out_0_11),
    .x                                                 (0),
    .y                                                 (11)
)vpe_0_11(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[0][11]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[0][11]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[0][11]),
    .cast_data_o                                       (cast_data_pe_2_nw[0][11]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[0][11]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[0][11]),
    .merge_data_i                                      (merge_data_nw_2_pe[0][11]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[0][11]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[0][11]),
    .merge_data_o                                      (merge_data_pe_2_nw[0][11]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[0][11]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[0][11]),
    .gather_data_i                                     (gather_data_nw_2_pe[0][11]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[0][11]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[0][11]),
    .gather_data_o                                     (gather_data_pe_2_nw[0][11]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[0][11]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[0][11])
);


virtual_pe #(
    .cast_out                                          (cast_out_0_12),
    .merge_in                                          (merge_in_0_12),
    .merge_out                                         (merge_out_0_12),
    .gather_in                                         (gather_in_0_12),
    .gather_out                                        (gather_out_0_12),
    .x                                                 (0),
    .y                                                 (12)
)vpe_0_12(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[0][12]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[0][12]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[0][12]),
    .cast_data_o                                       (cast_data_pe_2_nw[0][12]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[0][12]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[0][12]),
    .merge_data_i                                      (merge_data_nw_2_pe[0][12]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[0][12]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[0][12]),
    .merge_data_o                                      (merge_data_pe_2_nw[0][12]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[0][12]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[0][12]),
    .gather_data_i                                     (gather_data_nw_2_pe[0][12]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[0][12]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[0][12]),
    .gather_data_o                                     (gather_data_pe_2_nw[0][12]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[0][12]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[0][12])
);


virtual_pe #(
    .cast_out                                          (cast_out_0_13),
    .merge_in                                          (merge_in_0_13),
    .merge_out                                         (merge_out_0_13),
    .gather_in                                         (gather_in_0_13),
    .gather_out                                        (gather_out_0_13),
    .x                                                 (0),
    .y                                                 (13)
)vpe_0_13(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[0][13]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[0][13]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[0][13]),
    .cast_data_o                                       (cast_data_pe_2_nw[0][13]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[0][13]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[0][13]),
    .merge_data_i                                      (merge_data_nw_2_pe[0][13]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[0][13]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[0][13]),
    .merge_data_o                                      (merge_data_pe_2_nw[0][13]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[0][13]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[0][13]),
    .gather_data_i                                     (gather_data_nw_2_pe[0][13]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[0][13]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[0][13]),
    .gather_data_o                                     (gather_data_pe_2_nw[0][13]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[0][13]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[0][13])
);


virtual_pe #(
    .cast_out                                          (cast_out_0_14),
    .merge_in                                          (merge_in_0_14),
    .merge_out                                         (merge_out_0_14),
    .gather_in                                         (gather_in_0_14),
    .gather_out                                        (gather_out_0_14),
    .x                                                 (0),
    .y                                                 (14)
)vpe_0_14(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[0][14]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[0][14]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[0][14]),
    .cast_data_o                                       (cast_data_pe_2_nw[0][14]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[0][14]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[0][14]),
    .merge_data_i                                      (merge_data_nw_2_pe[0][14]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[0][14]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[0][14]),
    .merge_data_o                                      (merge_data_pe_2_nw[0][14]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[0][14]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[0][14]),
    .gather_data_i                                     (gather_data_nw_2_pe[0][14]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[0][14]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[0][14]),
    .gather_data_o                                     (gather_data_pe_2_nw[0][14]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[0][14]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[0][14])
);


virtual_pe #(
    .cast_out                                          (cast_out_0_15),
    .merge_in                                          (merge_in_0_15),
    .merge_out                                         (merge_out_0_15),
    .gather_in                                         (gather_in_0_15),
    .gather_out                                        (gather_out_0_15),
    .x                                                 (0),
    .y                                                 (15)
)vpe_0_15(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[0][15]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[0][15]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[0][15]),
    .cast_data_o                                       (cast_data_pe_2_nw[0][15]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[0][15]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[0][15]),
    .merge_data_i                                      (merge_data_nw_2_pe[0][15]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[0][15]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[0][15]),
    .merge_data_o                                      (merge_data_pe_2_nw[0][15]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[0][15]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[0][15]),
    .gather_data_i                                     (gather_data_nw_2_pe[0][15]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[0][15]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[0][15]),
    .gather_data_o                                     (gather_data_pe_2_nw[0][15]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[0][15]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[0][15])
);


virtual_pe #(
    .cast_out                                          (cast_out_0_16),
    .merge_in                                          (merge_in_0_16),
    .merge_out                                         (merge_out_0_16),
    .gather_in                                         (gather_in_0_16),
    .gather_out                                        (gather_out_0_16),
    .x                                                 (0),
    .y                                                 (16)
)vpe_0_16(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[0][16]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[0][16]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[0][16]),
    .cast_data_o                                       (cast_data_pe_2_nw[0][16]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[0][16]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[0][16]),
    .merge_data_i                                      (merge_data_nw_2_pe[0][16]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[0][16]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[0][16]),
    .merge_data_o                                      (merge_data_pe_2_nw[0][16]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[0][16]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[0][16]),
    .gather_data_i                                     (gather_data_nw_2_pe[0][16]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[0][16]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[0][16]),
    .gather_data_o                                     (gather_data_pe_2_nw[0][16]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[0][16]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[0][16])
);


virtual_pe #(
    .cast_out                                          (cast_out_0_17),
    .merge_in                                          (merge_in_0_17),
    .merge_out                                         (merge_out_0_17),
    .gather_in                                         (gather_in_0_17),
    .gather_out                                        (gather_out_0_17),
    .x                                                 (0),
    .y                                                 (17)
)vpe_0_17(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[0][17]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[0][17]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[0][17]),
    .cast_data_o                                       (cast_data_pe_2_nw[0][17]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[0][17]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[0][17]),
    .merge_data_i                                      (merge_data_nw_2_pe[0][17]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[0][17]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[0][17]),
    .merge_data_o                                      (merge_data_pe_2_nw[0][17]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[0][17]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[0][17]),
    .gather_data_i                                     (gather_data_nw_2_pe[0][17]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[0][17]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[0][17]),
    .gather_data_o                                     (gather_data_pe_2_nw[0][17]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[0][17]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[0][17])
);


virtual_pe #(
    .cast_out                                          (cast_out_0_18),
    .merge_in                                          (merge_in_0_18),
    .merge_out                                         (merge_out_0_18),
    .gather_in                                         (gather_in_0_18),
    .gather_out                                        (gather_out_0_18),
    .x                                                 (0),
    .y                                                 (18)
)vpe_0_18(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[0][18]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[0][18]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[0][18]),
    .cast_data_o                                       (cast_data_pe_2_nw[0][18]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[0][18]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[0][18]),
    .merge_data_i                                      (merge_data_nw_2_pe[0][18]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[0][18]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[0][18]),
    .merge_data_o                                      (merge_data_pe_2_nw[0][18]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[0][18]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[0][18]),
    .gather_data_i                                     (gather_data_nw_2_pe[0][18]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[0][18]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[0][18]),
    .gather_data_o                                     (gather_data_pe_2_nw[0][18]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[0][18]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[0][18])
);


virtual_pe #(
    .cast_out                                          (cast_out_0_19),
    .merge_in                                          (merge_in_0_19),
    .merge_out                                         (merge_out_0_19),
    .gather_in                                         (gather_in_0_19),
    .gather_out                                        (gather_out_0_19),
    .x                                                 (0),
    .y                                                 (19)
)vpe_0_19(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[0][19]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[0][19]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[0][19]),
    .cast_data_o                                       (cast_data_pe_2_nw[0][19]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[0][19]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[0][19]),
    .merge_data_i                                      (merge_data_nw_2_pe[0][19]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[0][19]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[0][19]),
    .merge_data_o                                      (merge_data_pe_2_nw[0][19]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[0][19]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[0][19]),
    .gather_data_i                                     (gather_data_nw_2_pe[0][19]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[0][19]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[0][19]),
    .gather_data_o                                     (gather_data_pe_2_nw[0][19]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[0][19]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[0][19])
);


virtual_pe #(
    .cast_out                                          (cast_out_0_20),
    .merge_in                                          (merge_in_0_20),
    .merge_out                                         (merge_out_0_20),
    .gather_in                                         (gather_in_0_20),
    .gather_out                                        (gather_out_0_20),
    .x                                                 (0),
    .y                                                 (20)
)vpe_0_20(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[0][20]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[0][20]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[0][20]),
    .cast_data_o                                       (cast_data_pe_2_nw[0][20]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[0][20]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[0][20]),
    .merge_data_i                                      (merge_data_nw_2_pe[0][20]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[0][20]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[0][20]),
    .merge_data_o                                      (merge_data_pe_2_nw[0][20]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[0][20]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[0][20]),
    .gather_data_i                                     (gather_data_nw_2_pe[0][20]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[0][20]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[0][20]),
    .gather_data_o                                     (gather_data_pe_2_nw[0][20]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[0][20]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[0][20])
);


virtual_pe #(
    .cast_out                                          (cast_out_0_21),
    .merge_in                                          (merge_in_0_21),
    .merge_out                                         (merge_out_0_21),
    .gather_in                                         (gather_in_0_21),
    .gather_out                                        (gather_out_0_21),
    .x                                                 (0),
    .y                                                 (21)
)vpe_0_21(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[0][21]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[0][21]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[0][21]),
    .cast_data_o                                       (cast_data_pe_2_nw[0][21]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[0][21]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[0][21]),
    .merge_data_i                                      (merge_data_nw_2_pe[0][21]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[0][21]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[0][21]),
    .merge_data_o                                      (merge_data_pe_2_nw[0][21]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[0][21]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[0][21]),
    .gather_data_i                                     (gather_data_nw_2_pe[0][21]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[0][21]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[0][21]),
    .gather_data_o                                     (gather_data_pe_2_nw[0][21]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[0][21]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[0][21])
);


virtual_pe #(
    .cast_out                                          (cast_out_0_22),
    .merge_in                                          (merge_in_0_22),
    .merge_out                                         (merge_out_0_22),
    .gather_in                                         (gather_in_0_22),
    .gather_out                                        (gather_out_0_22),
    .x                                                 (0),
    .y                                                 (22)
)vpe_0_22(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[0][22]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[0][22]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[0][22]),
    .cast_data_o                                       (cast_data_pe_2_nw[0][22]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[0][22]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[0][22]),
    .merge_data_i                                      (merge_data_nw_2_pe[0][22]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[0][22]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[0][22]),
    .merge_data_o                                      (merge_data_pe_2_nw[0][22]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[0][22]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[0][22]),
    .gather_data_i                                     (gather_data_nw_2_pe[0][22]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[0][22]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[0][22]),
    .gather_data_o                                     (gather_data_pe_2_nw[0][22]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[0][22]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[0][22])
);


virtual_pe #(
    .cast_out                                          (cast_out_0_23),
    .merge_in                                          (merge_in_0_23),
    .merge_out                                         (merge_out_0_23),
    .gather_in                                         (gather_in_0_23),
    .gather_out                                        (gather_out_0_23),
    .x                                                 (0),
    .y                                                 (23)
)vpe_0_23(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[0][23]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[0][23]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[0][23]),
    .cast_data_o                                       (cast_data_pe_2_nw[0][23]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[0][23]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[0][23]),
    .merge_data_i                                      (merge_data_nw_2_pe[0][23]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[0][23]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[0][23]),
    .merge_data_o                                      (merge_data_pe_2_nw[0][23]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[0][23]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[0][23]),
    .gather_data_i                                     (gather_data_nw_2_pe[0][23]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[0][23]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[0][23]),
    .gather_data_o                                     (gather_data_pe_2_nw[0][23]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[0][23]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[0][23])
);


virtual_pe #(
    .cast_out                                          (cast_out_0_24),
    .merge_in                                          (merge_in_0_24),
    .merge_out                                         (merge_out_0_24),
    .gather_in                                         (gather_in_0_24),
    .gather_out                                        (gather_out_0_24),
    .x                                                 (0),
    .y                                                 (24)
)vpe_0_24(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[0][24]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[0][24]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[0][24]),
    .cast_data_o                                       (cast_data_pe_2_nw[0][24]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[0][24]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[0][24]),
    .merge_data_i                                      (merge_data_nw_2_pe[0][24]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[0][24]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[0][24]),
    .merge_data_o                                      (merge_data_pe_2_nw[0][24]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[0][24]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[0][24]),
    .gather_data_i                                     (gather_data_nw_2_pe[0][24]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[0][24]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[0][24]),
    .gather_data_o                                     (gather_data_pe_2_nw[0][24]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[0][24]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[0][24])
);


virtual_pe #(
    .cast_out                                          (cast_out_1_0),
    .merge_in                                          (merge_in_1_0),
    .merge_out                                         (merge_out_1_0),
    .gather_in                                         (gather_in_1_0),
    .gather_out                                        (gather_out_1_0),
    .x                                                 (1),
    .y                                                 (0)
)vpe_1_0(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[1][0]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[1][0]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[1][0]),
    .cast_data_o                                       (cast_data_pe_2_nw[1][0]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[1][0]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[1][0]),
    .merge_data_i                                      (merge_data_nw_2_pe[1][0]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[1][0]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[1][0]),
    .merge_data_o                                      (merge_data_pe_2_nw[1][0]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[1][0]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[1][0]),
    .gather_data_i                                     (gather_data_nw_2_pe[1][0]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[1][0]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[1][0]),
    .gather_data_o                                     (gather_data_pe_2_nw[1][0]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[1][0]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[1][0])
);


virtual_pe #(
    .cast_out                                          (cast_out_1_1),
    .merge_in                                          (merge_in_1_1),
    .merge_out                                         (merge_out_1_1),
    .gather_in                                         (gather_in_1_1),
    .gather_out                                        (gather_out_1_1),
    .x                                                 (1),
    .y                                                 (1)
)vpe_1_1(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[1][1]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[1][1]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[1][1]),
    .cast_data_o                                       (cast_data_pe_2_nw[1][1]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[1][1]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[1][1]),
    .merge_data_i                                      (merge_data_nw_2_pe[1][1]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[1][1]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[1][1]),
    .merge_data_o                                      (merge_data_pe_2_nw[1][1]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[1][1]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[1][1]),
    .gather_data_i                                     (gather_data_nw_2_pe[1][1]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[1][1]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[1][1]),
    .gather_data_o                                     (gather_data_pe_2_nw[1][1]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[1][1]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[1][1])
);


virtual_pe #(
    .cast_out                                          (cast_out_1_2),
    .merge_in                                          (merge_in_1_2),
    .merge_out                                         (merge_out_1_2),
    .gather_in                                         (gather_in_1_2),
    .gather_out                                        (gather_out_1_2),
    .x                                                 (1),
    .y                                                 (2)
)vpe_1_2(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[1][2]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[1][2]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[1][2]),
    .cast_data_o                                       (cast_data_pe_2_nw[1][2]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[1][2]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[1][2]),
    .merge_data_i                                      (merge_data_nw_2_pe[1][2]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[1][2]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[1][2]),
    .merge_data_o                                      (merge_data_pe_2_nw[1][2]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[1][2]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[1][2]),
    .gather_data_i                                     (gather_data_nw_2_pe[1][2]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[1][2]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[1][2]),
    .gather_data_o                                     (gather_data_pe_2_nw[1][2]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[1][2]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[1][2])
);


virtual_pe #(
    .cast_out                                          (cast_out_1_3),
    .merge_in                                          (merge_in_1_3),
    .merge_out                                         (merge_out_1_3),
    .gather_in                                         (gather_in_1_3),
    .gather_out                                        (gather_out_1_3),
    .x                                                 (1),
    .y                                                 (3)
)vpe_1_3(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[1][3]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[1][3]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[1][3]),
    .cast_data_o                                       (cast_data_pe_2_nw[1][3]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[1][3]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[1][3]),
    .merge_data_i                                      (merge_data_nw_2_pe[1][3]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[1][3]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[1][3]),
    .merge_data_o                                      (merge_data_pe_2_nw[1][3]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[1][3]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[1][3]),
    .gather_data_i                                     (gather_data_nw_2_pe[1][3]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[1][3]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[1][3]),
    .gather_data_o                                     (gather_data_pe_2_nw[1][3]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[1][3]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[1][3])
);


virtual_pe #(
    .cast_out                                          (cast_out_1_4),
    .merge_in                                          (merge_in_1_4),
    .merge_out                                         (merge_out_1_4),
    .gather_in                                         (gather_in_1_4),
    .gather_out                                        (gather_out_1_4),
    .x                                                 (1),
    .y                                                 (4)
)vpe_1_4(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[1][4]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[1][4]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[1][4]),
    .cast_data_o                                       (cast_data_pe_2_nw[1][4]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[1][4]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[1][4]),
    .merge_data_i                                      (merge_data_nw_2_pe[1][4]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[1][4]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[1][4]),
    .merge_data_o                                      (merge_data_pe_2_nw[1][4]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[1][4]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[1][4]),
    .gather_data_i                                     (gather_data_nw_2_pe[1][4]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[1][4]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[1][4]),
    .gather_data_o                                     (gather_data_pe_2_nw[1][4]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[1][4]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[1][4])
);


virtual_pe #(
    .cast_out                                          (cast_out_1_5),
    .merge_in                                          (merge_in_1_5),
    .merge_out                                         (merge_out_1_5),
    .gather_in                                         (gather_in_1_5),
    .gather_out                                        (gather_out_1_5),
    .x                                                 (1),
    .y                                                 (5)
)vpe_1_5(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[1][5]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[1][5]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[1][5]),
    .cast_data_o                                       (cast_data_pe_2_nw[1][5]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[1][5]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[1][5]),
    .merge_data_i                                      (merge_data_nw_2_pe[1][5]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[1][5]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[1][5]),
    .merge_data_o                                      (merge_data_pe_2_nw[1][5]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[1][5]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[1][5]),
    .gather_data_i                                     (gather_data_nw_2_pe[1][5]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[1][5]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[1][5]),
    .gather_data_o                                     (gather_data_pe_2_nw[1][5]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[1][5]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[1][5])
);


virtual_pe #(
    .cast_out                                          (cast_out_1_6),
    .merge_in                                          (merge_in_1_6),
    .merge_out                                         (merge_out_1_6),
    .gather_in                                         (gather_in_1_6),
    .gather_out                                        (gather_out_1_6),
    .x                                                 (1),
    .y                                                 (6)
)vpe_1_6(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[1][6]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[1][6]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[1][6]),
    .cast_data_o                                       (cast_data_pe_2_nw[1][6]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[1][6]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[1][6]),
    .merge_data_i                                      (merge_data_nw_2_pe[1][6]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[1][6]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[1][6]),
    .merge_data_o                                      (merge_data_pe_2_nw[1][6]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[1][6]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[1][6]),
    .gather_data_i                                     (gather_data_nw_2_pe[1][6]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[1][6]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[1][6]),
    .gather_data_o                                     (gather_data_pe_2_nw[1][6]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[1][6]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[1][6])
);


virtual_pe #(
    .cast_out                                          (cast_out_1_7),
    .merge_in                                          (merge_in_1_7),
    .merge_out                                         (merge_out_1_7),
    .gather_in                                         (gather_in_1_7),
    .gather_out                                        (gather_out_1_7),
    .x                                                 (1),
    .y                                                 (7)
)vpe_1_7(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[1][7]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[1][7]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[1][7]),
    .cast_data_o                                       (cast_data_pe_2_nw[1][7]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[1][7]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[1][7]),
    .merge_data_i                                      (merge_data_nw_2_pe[1][7]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[1][7]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[1][7]),
    .merge_data_o                                      (merge_data_pe_2_nw[1][7]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[1][7]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[1][7]),
    .gather_data_i                                     (gather_data_nw_2_pe[1][7]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[1][7]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[1][7]),
    .gather_data_o                                     (gather_data_pe_2_nw[1][7]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[1][7]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[1][7])
);


virtual_pe #(
    .cast_out                                          (cast_out_1_8),
    .merge_in                                          (merge_in_1_8),
    .merge_out                                         (merge_out_1_8),
    .gather_in                                         (gather_in_1_8),
    .gather_out                                        (gather_out_1_8),
    .x                                                 (1),
    .y                                                 (8)
)vpe_1_8(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[1][8]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[1][8]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[1][8]),
    .cast_data_o                                       (cast_data_pe_2_nw[1][8]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[1][8]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[1][8]),
    .merge_data_i                                      (merge_data_nw_2_pe[1][8]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[1][8]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[1][8]),
    .merge_data_o                                      (merge_data_pe_2_nw[1][8]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[1][8]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[1][8]),
    .gather_data_i                                     (gather_data_nw_2_pe[1][8]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[1][8]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[1][8]),
    .gather_data_o                                     (gather_data_pe_2_nw[1][8]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[1][8]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[1][8])
);


virtual_pe #(
    .cast_out                                          (cast_out_1_9),
    .merge_in                                          (merge_in_1_9),
    .merge_out                                         (merge_out_1_9),
    .gather_in                                         (gather_in_1_9),
    .gather_out                                        (gather_out_1_9),
    .x                                                 (1),
    .y                                                 (9)
)vpe_1_9(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[1][9]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[1][9]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[1][9]),
    .cast_data_o                                       (cast_data_pe_2_nw[1][9]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[1][9]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[1][9]),
    .merge_data_i                                      (merge_data_nw_2_pe[1][9]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[1][9]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[1][9]),
    .merge_data_o                                      (merge_data_pe_2_nw[1][9]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[1][9]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[1][9]),
    .gather_data_i                                     (gather_data_nw_2_pe[1][9]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[1][9]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[1][9]),
    .gather_data_o                                     (gather_data_pe_2_nw[1][9]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[1][9]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[1][9])
);


virtual_pe #(
    .cast_out                                          (cast_out_1_10),
    .merge_in                                          (merge_in_1_10),
    .merge_out                                         (merge_out_1_10),
    .gather_in                                         (gather_in_1_10),
    .gather_out                                        (gather_out_1_10),
    .x                                                 (1),
    .y                                                 (10)
)vpe_1_10(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[1][10]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[1][10]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[1][10]),
    .cast_data_o                                       (cast_data_pe_2_nw[1][10]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[1][10]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[1][10]),
    .merge_data_i                                      (merge_data_nw_2_pe[1][10]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[1][10]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[1][10]),
    .merge_data_o                                      (merge_data_pe_2_nw[1][10]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[1][10]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[1][10]),
    .gather_data_i                                     (gather_data_nw_2_pe[1][10]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[1][10]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[1][10]),
    .gather_data_o                                     (gather_data_pe_2_nw[1][10]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[1][10]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[1][10])
);


virtual_pe #(
    .cast_out                                          (cast_out_1_11),
    .merge_in                                          (merge_in_1_11),
    .merge_out                                         (merge_out_1_11),
    .gather_in                                         (gather_in_1_11),
    .gather_out                                        (gather_out_1_11),
    .x                                                 (1),
    .y                                                 (11)
)vpe_1_11(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[1][11]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[1][11]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[1][11]),
    .cast_data_o                                       (cast_data_pe_2_nw[1][11]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[1][11]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[1][11]),
    .merge_data_i                                      (merge_data_nw_2_pe[1][11]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[1][11]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[1][11]),
    .merge_data_o                                      (merge_data_pe_2_nw[1][11]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[1][11]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[1][11]),
    .gather_data_i                                     (gather_data_nw_2_pe[1][11]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[1][11]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[1][11]),
    .gather_data_o                                     (gather_data_pe_2_nw[1][11]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[1][11]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[1][11])
);


virtual_pe #(
    .cast_out                                          (cast_out_1_12),
    .merge_in                                          (merge_in_1_12),
    .merge_out                                         (merge_out_1_12),
    .gather_in                                         (gather_in_1_12),
    .gather_out                                        (gather_out_1_12),
    .x                                                 (1),
    .y                                                 (12)
)vpe_1_12(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[1][12]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[1][12]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[1][12]),
    .cast_data_o                                       (cast_data_pe_2_nw[1][12]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[1][12]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[1][12]),
    .merge_data_i                                      (merge_data_nw_2_pe[1][12]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[1][12]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[1][12]),
    .merge_data_o                                      (merge_data_pe_2_nw[1][12]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[1][12]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[1][12]),
    .gather_data_i                                     (gather_data_nw_2_pe[1][12]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[1][12]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[1][12]),
    .gather_data_o                                     (gather_data_pe_2_nw[1][12]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[1][12]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[1][12])
);


virtual_pe #(
    .cast_out                                          (cast_out_1_13),
    .merge_in                                          (merge_in_1_13),
    .merge_out                                         (merge_out_1_13),
    .gather_in                                         (gather_in_1_13),
    .gather_out                                        (gather_out_1_13),
    .x                                                 (1),
    .y                                                 (13)
)vpe_1_13(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[1][13]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[1][13]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[1][13]),
    .cast_data_o                                       (cast_data_pe_2_nw[1][13]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[1][13]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[1][13]),
    .merge_data_i                                      (merge_data_nw_2_pe[1][13]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[1][13]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[1][13]),
    .merge_data_o                                      (merge_data_pe_2_nw[1][13]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[1][13]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[1][13]),
    .gather_data_i                                     (gather_data_nw_2_pe[1][13]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[1][13]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[1][13]),
    .gather_data_o                                     (gather_data_pe_2_nw[1][13]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[1][13]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[1][13])
);


virtual_pe #(
    .cast_out                                          (cast_out_1_14),
    .merge_in                                          (merge_in_1_14),
    .merge_out                                         (merge_out_1_14),
    .gather_in                                         (gather_in_1_14),
    .gather_out                                        (gather_out_1_14),
    .x                                                 (1),
    .y                                                 (14)
)vpe_1_14(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[1][14]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[1][14]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[1][14]),
    .cast_data_o                                       (cast_data_pe_2_nw[1][14]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[1][14]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[1][14]),
    .merge_data_i                                      (merge_data_nw_2_pe[1][14]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[1][14]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[1][14]),
    .merge_data_o                                      (merge_data_pe_2_nw[1][14]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[1][14]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[1][14]),
    .gather_data_i                                     (gather_data_nw_2_pe[1][14]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[1][14]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[1][14]),
    .gather_data_o                                     (gather_data_pe_2_nw[1][14]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[1][14]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[1][14])
);


virtual_pe #(
    .cast_out                                          (cast_out_1_15),
    .merge_in                                          (merge_in_1_15),
    .merge_out                                         (merge_out_1_15),
    .gather_in                                         (gather_in_1_15),
    .gather_out                                        (gather_out_1_15),
    .x                                                 (1),
    .y                                                 (15)
)vpe_1_15(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[1][15]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[1][15]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[1][15]),
    .cast_data_o                                       (cast_data_pe_2_nw[1][15]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[1][15]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[1][15]),
    .merge_data_i                                      (merge_data_nw_2_pe[1][15]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[1][15]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[1][15]),
    .merge_data_o                                      (merge_data_pe_2_nw[1][15]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[1][15]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[1][15]),
    .gather_data_i                                     (gather_data_nw_2_pe[1][15]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[1][15]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[1][15]),
    .gather_data_o                                     (gather_data_pe_2_nw[1][15]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[1][15]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[1][15])
);


virtual_pe #(
    .cast_out                                          (cast_out_1_16),
    .merge_in                                          (merge_in_1_16),
    .merge_out                                         (merge_out_1_16),
    .gather_in                                         (gather_in_1_16),
    .gather_out                                        (gather_out_1_16),
    .x                                                 (1),
    .y                                                 (16)
)vpe_1_16(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[1][16]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[1][16]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[1][16]),
    .cast_data_o                                       (cast_data_pe_2_nw[1][16]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[1][16]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[1][16]),
    .merge_data_i                                      (merge_data_nw_2_pe[1][16]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[1][16]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[1][16]),
    .merge_data_o                                      (merge_data_pe_2_nw[1][16]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[1][16]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[1][16]),
    .gather_data_i                                     (gather_data_nw_2_pe[1][16]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[1][16]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[1][16]),
    .gather_data_o                                     (gather_data_pe_2_nw[1][16]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[1][16]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[1][16])
);


virtual_pe #(
    .cast_out                                          (cast_out_1_17),
    .merge_in                                          (merge_in_1_17),
    .merge_out                                         (merge_out_1_17),
    .gather_in                                         (gather_in_1_17),
    .gather_out                                        (gather_out_1_17),
    .x                                                 (1),
    .y                                                 (17)
)vpe_1_17(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[1][17]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[1][17]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[1][17]),
    .cast_data_o                                       (cast_data_pe_2_nw[1][17]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[1][17]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[1][17]),
    .merge_data_i                                      (merge_data_nw_2_pe[1][17]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[1][17]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[1][17]),
    .merge_data_o                                      (merge_data_pe_2_nw[1][17]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[1][17]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[1][17]),
    .gather_data_i                                     (gather_data_nw_2_pe[1][17]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[1][17]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[1][17]),
    .gather_data_o                                     (gather_data_pe_2_nw[1][17]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[1][17]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[1][17])
);


virtual_pe #(
    .cast_out                                          (cast_out_1_18),
    .merge_in                                          (merge_in_1_18),
    .merge_out                                         (merge_out_1_18),
    .gather_in                                         (gather_in_1_18),
    .gather_out                                        (gather_out_1_18),
    .x                                                 (1),
    .y                                                 (18)
)vpe_1_18(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[1][18]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[1][18]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[1][18]),
    .cast_data_o                                       (cast_data_pe_2_nw[1][18]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[1][18]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[1][18]),
    .merge_data_i                                      (merge_data_nw_2_pe[1][18]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[1][18]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[1][18]),
    .merge_data_o                                      (merge_data_pe_2_nw[1][18]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[1][18]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[1][18]),
    .gather_data_i                                     (gather_data_nw_2_pe[1][18]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[1][18]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[1][18]),
    .gather_data_o                                     (gather_data_pe_2_nw[1][18]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[1][18]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[1][18])
);


virtual_pe #(
    .cast_out                                          (cast_out_1_19),
    .merge_in                                          (merge_in_1_19),
    .merge_out                                         (merge_out_1_19),
    .gather_in                                         (gather_in_1_19),
    .gather_out                                        (gather_out_1_19),
    .x                                                 (1),
    .y                                                 (19)
)vpe_1_19(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[1][19]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[1][19]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[1][19]),
    .cast_data_o                                       (cast_data_pe_2_nw[1][19]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[1][19]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[1][19]),
    .merge_data_i                                      (merge_data_nw_2_pe[1][19]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[1][19]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[1][19]),
    .merge_data_o                                      (merge_data_pe_2_nw[1][19]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[1][19]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[1][19]),
    .gather_data_i                                     (gather_data_nw_2_pe[1][19]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[1][19]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[1][19]),
    .gather_data_o                                     (gather_data_pe_2_nw[1][19]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[1][19]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[1][19])
);


virtual_pe #(
    .cast_out                                          (cast_out_1_20),
    .merge_in                                          (merge_in_1_20),
    .merge_out                                         (merge_out_1_20),
    .gather_in                                         (gather_in_1_20),
    .gather_out                                        (gather_out_1_20),
    .x                                                 (1),
    .y                                                 (20)
)vpe_1_20(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[1][20]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[1][20]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[1][20]),
    .cast_data_o                                       (cast_data_pe_2_nw[1][20]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[1][20]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[1][20]),
    .merge_data_i                                      (merge_data_nw_2_pe[1][20]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[1][20]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[1][20]),
    .merge_data_o                                      (merge_data_pe_2_nw[1][20]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[1][20]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[1][20]),
    .gather_data_i                                     (gather_data_nw_2_pe[1][20]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[1][20]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[1][20]),
    .gather_data_o                                     (gather_data_pe_2_nw[1][20]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[1][20]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[1][20])
);


virtual_pe #(
    .cast_out                                          (cast_out_1_21),
    .merge_in                                          (merge_in_1_21),
    .merge_out                                         (merge_out_1_21),
    .gather_in                                         (gather_in_1_21),
    .gather_out                                        (gather_out_1_21),
    .x                                                 (1),
    .y                                                 (21)
)vpe_1_21(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[1][21]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[1][21]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[1][21]),
    .cast_data_o                                       (cast_data_pe_2_nw[1][21]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[1][21]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[1][21]),
    .merge_data_i                                      (merge_data_nw_2_pe[1][21]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[1][21]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[1][21]),
    .merge_data_o                                      (merge_data_pe_2_nw[1][21]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[1][21]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[1][21]),
    .gather_data_i                                     (gather_data_nw_2_pe[1][21]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[1][21]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[1][21]),
    .gather_data_o                                     (gather_data_pe_2_nw[1][21]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[1][21]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[1][21])
);


virtual_pe #(
    .cast_out                                          (cast_out_1_22),
    .merge_in                                          (merge_in_1_22),
    .merge_out                                         (merge_out_1_22),
    .gather_in                                         (gather_in_1_22),
    .gather_out                                        (gather_out_1_22),
    .x                                                 (1),
    .y                                                 (22)
)vpe_1_22(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[1][22]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[1][22]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[1][22]),
    .cast_data_o                                       (cast_data_pe_2_nw[1][22]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[1][22]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[1][22]),
    .merge_data_i                                      (merge_data_nw_2_pe[1][22]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[1][22]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[1][22]),
    .merge_data_o                                      (merge_data_pe_2_nw[1][22]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[1][22]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[1][22]),
    .gather_data_i                                     (gather_data_nw_2_pe[1][22]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[1][22]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[1][22]),
    .gather_data_o                                     (gather_data_pe_2_nw[1][22]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[1][22]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[1][22])
);


virtual_pe #(
    .cast_out                                          (cast_out_1_23),
    .merge_in                                          (merge_in_1_23),
    .merge_out                                         (merge_out_1_23),
    .gather_in                                         (gather_in_1_23),
    .gather_out                                        (gather_out_1_23),
    .x                                                 (1),
    .y                                                 (23)
)vpe_1_23(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[1][23]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[1][23]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[1][23]),
    .cast_data_o                                       (cast_data_pe_2_nw[1][23]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[1][23]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[1][23]),
    .merge_data_i                                      (merge_data_nw_2_pe[1][23]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[1][23]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[1][23]),
    .merge_data_o                                      (merge_data_pe_2_nw[1][23]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[1][23]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[1][23]),
    .gather_data_i                                     (gather_data_nw_2_pe[1][23]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[1][23]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[1][23]),
    .gather_data_o                                     (gather_data_pe_2_nw[1][23]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[1][23]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[1][23])
);


virtual_pe #(
    .cast_out                                          (cast_out_1_24),
    .merge_in                                          (merge_in_1_24),
    .merge_out                                         (merge_out_1_24),
    .gather_in                                         (gather_in_1_24),
    .gather_out                                        (gather_out_1_24),
    .x                                                 (1),
    .y                                                 (24)
)vpe_1_24(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[1][24]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[1][24]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[1][24]),
    .cast_data_o                                       (cast_data_pe_2_nw[1][24]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[1][24]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[1][24]),
    .merge_data_i                                      (merge_data_nw_2_pe[1][24]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[1][24]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[1][24]),
    .merge_data_o                                      (merge_data_pe_2_nw[1][24]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[1][24]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[1][24]),
    .gather_data_i                                     (gather_data_nw_2_pe[1][24]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[1][24]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[1][24]),
    .gather_data_o                                     (gather_data_pe_2_nw[1][24]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[1][24]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[1][24])
);


virtual_pe #(
    .cast_out                                          (cast_out_2_0),
    .merge_in                                          (merge_in_2_0),
    .merge_out                                         (merge_out_2_0),
    .gather_in                                         (gather_in_2_0),
    .gather_out                                        (gather_out_2_0),
    .x                                                 (2),
    .y                                                 (0)
)vpe_2_0(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[2][0]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[2][0]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[2][0]),
    .cast_data_o                                       (cast_data_pe_2_nw[2][0]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[2][0]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[2][0]),
    .merge_data_i                                      (merge_data_nw_2_pe[2][0]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[2][0]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[2][0]),
    .merge_data_o                                      (merge_data_pe_2_nw[2][0]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[2][0]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[2][0]),
    .gather_data_i                                     (gather_data_nw_2_pe[2][0]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[2][0]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[2][0]),
    .gather_data_o                                     (gather_data_pe_2_nw[2][0]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[2][0]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[2][0])
);


virtual_pe #(
    .cast_out                                          (cast_out_2_1),
    .merge_in                                          (merge_in_2_1),
    .merge_out                                         (merge_out_2_1),
    .gather_in                                         (gather_in_2_1),
    .gather_out                                        (gather_out_2_1),
    .x                                                 (2),
    .y                                                 (1)
)vpe_2_1(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[2][1]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[2][1]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[2][1]),
    .cast_data_o                                       (cast_data_pe_2_nw[2][1]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[2][1]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[2][1]),
    .merge_data_i                                      (merge_data_nw_2_pe[2][1]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[2][1]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[2][1]),
    .merge_data_o                                      (merge_data_pe_2_nw[2][1]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[2][1]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[2][1]),
    .gather_data_i                                     (gather_data_nw_2_pe[2][1]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[2][1]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[2][1]),
    .gather_data_o                                     (gather_data_pe_2_nw[2][1]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[2][1]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[2][1])
);


virtual_pe #(
    .cast_out                                          (cast_out_2_2),
    .merge_in                                          (merge_in_2_2),
    .merge_out                                         (merge_out_2_2),
    .gather_in                                         (gather_in_2_2),
    .gather_out                                        (gather_out_2_2),
    .x                                                 (2),
    .y                                                 (2)
)vpe_2_2(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[2][2]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[2][2]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[2][2]),
    .cast_data_o                                       (cast_data_pe_2_nw[2][2]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[2][2]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[2][2]),
    .merge_data_i                                      (merge_data_nw_2_pe[2][2]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[2][2]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[2][2]),
    .merge_data_o                                      (merge_data_pe_2_nw[2][2]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[2][2]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[2][2]),
    .gather_data_i                                     (gather_data_nw_2_pe[2][2]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[2][2]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[2][2]),
    .gather_data_o                                     (gather_data_pe_2_nw[2][2]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[2][2]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[2][2])
);


virtual_pe #(
    .cast_out                                          (cast_out_2_3),
    .merge_in                                          (merge_in_2_3),
    .merge_out                                         (merge_out_2_3),
    .gather_in                                         (gather_in_2_3),
    .gather_out                                        (gather_out_2_3),
    .x                                                 (2),
    .y                                                 (3)
)vpe_2_3(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[2][3]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[2][3]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[2][3]),
    .cast_data_o                                       (cast_data_pe_2_nw[2][3]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[2][3]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[2][3]),
    .merge_data_i                                      (merge_data_nw_2_pe[2][3]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[2][3]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[2][3]),
    .merge_data_o                                      (merge_data_pe_2_nw[2][3]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[2][3]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[2][3]),
    .gather_data_i                                     (gather_data_nw_2_pe[2][3]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[2][3]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[2][3]),
    .gather_data_o                                     (gather_data_pe_2_nw[2][3]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[2][3]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[2][3])
);


virtual_pe #(
    .cast_out                                          (cast_out_2_4),
    .merge_in                                          (merge_in_2_4),
    .merge_out                                         (merge_out_2_4),
    .gather_in                                         (gather_in_2_4),
    .gather_out                                        (gather_out_2_4),
    .x                                                 (2),
    .y                                                 (4)
)vpe_2_4(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[2][4]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[2][4]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[2][4]),
    .cast_data_o                                       (cast_data_pe_2_nw[2][4]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[2][4]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[2][4]),
    .merge_data_i                                      (merge_data_nw_2_pe[2][4]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[2][4]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[2][4]),
    .merge_data_o                                      (merge_data_pe_2_nw[2][4]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[2][4]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[2][4]),
    .gather_data_i                                     (gather_data_nw_2_pe[2][4]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[2][4]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[2][4]),
    .gather_data_o                                     (gather_data_pe_2_nw[2][4]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[2][4]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[2][4])
);


virtual_pe #(
    .cast_out                                          (cast_out_2_5),
    .merge_in                                          (merge_in_2_5),
    .merge_out                                         (merge_out_2_5),
    .gather_in                                         (gather_in_2_5),
    .gather_out                                        (gather_out_2_5),
    .x                                                 (2),
    .y                                                 (5)
)vpe_2_5(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[2][5]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[2][5]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[2][5]),
    .cast_data_o                                       (cast_data_pe_2_nw[2][5]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[2][5]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[2][5]),
    .merge_data_i                                      (merge_data_nw_2_pe[2][5]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[2][5]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[2][5]),
    .merge_data_o                                      (merge_data_pe_2_nw[2][5]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[2][5]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[2][5]),
    .gather_data_i                                     (gather_data_nw_2_pe[2][5]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[2][5]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[2][5]),
    .gather_data_o                                     (gather_data_pe_2_nw[2][5]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[2][5]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[2][5])
);


virtual_pe #(
    .cast_out                                          (cast_out_2_6),
    .merge_in                                          (merge_in_2_6),
    .merge_out                                         (merge_out_2_6),
    .gather_in                                         (gather_in_2_6),
    .gather_out                                        (gather_out_2_6),
    .x                                                 (2),
    .y                                                 (6)
)vpe_2_6(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[2][6]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[2][6]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[2][6]),
    .cast_data_o                                       (cast_data_pe_2_nw[2][6]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[2][6]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[2][6]),
    .merge_data_i                                      (merge_data_nw_2_pe[2][6]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[2][6]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[2][6]),
    .merge_data_o                                      (merge_data_pe_2_nw[2][6]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[2][6]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[2][6]),
    .gather_data_i                                     (gather_data_nw_2_pe[2][6]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[2][6]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[2][6]),
    .gather_data_o                                     (gather_data_pe_2_nw[2][6]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[2][6]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[2][6])
);


virtual_pe #(
    .cast_out                                          (cast_out_2_7),
    .merge_in                                          (merge_in_2_7),
    .merge_out                                         (merge_out_2_7),
    .gather_in                                         (gather_in_2_7),
    .gather_out                                        (gather_out_2_7),
    .x                                                 (2),
    .y                                                 (7)
)vpe_2_7(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[2][7]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[2][7]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[2][7]),
    .cast_data_o                                       (cast_data_pe_2_nw[2][7]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[2][7]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[2][7]),
    .merge_data_i                                      (merge_data_nw_2_pe[2][7]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[2][7]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[2][7]),
    .merge_data_o                                      (merge_data_pe_2_nw[2][7]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[2][7]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[2][7]),
    .gather_data_i                                     (gather_data_nw_2_pe[2][7]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[2][7]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[2][7]),
    .gather_data_o                                     (gather_data_pe_2_nw[2][7]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[2][7]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[2][7])
);


virtual_pe #(
    .cast_out                                          (cast_out_2_8),
    .merge_in                                          (merge_in_2_8),
    .merge_out                                         (merge_out_2_8),
    .gather_in                                         (gather_in_2_8),
    .gather_out                                        (gather_out_2_8),
    .x                                                 (2),
    .y                                                 (8)
)vpe_2_8(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[2][8]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[2][8]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[2][8]),
    .cast_data_o                                       (cast_data_pe_2_nw[2][8]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[2][8]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[2][8]),
    .merge_data_i                                      (merge_data_nw_2_pe[2][8]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[2][8]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[2][8]),
    .merge_data_o                                      (merge_data_pe_2_nw[2][8]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[2][8]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[2][8]),
    .gather_data_i                                     (gather_data_nw_2_pe[2][8]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[2][8]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[2][8]),
    .gather_data_o                                     (gather_data_pe_2_nw[2][8]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[2][8]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[2][8])
);


virtual_pe #(
    .cast_out                                          (cast_out_2_9),
    .merge_in                                          (merge_in_2_9),
    .merge_out                                         (merge_out_2_9),
    .gather_in                                         (gather_in_2_9),
    .gather_out                                        (gather_out_2_9),
    .x                                                 (2),
    .y                                                 (9)
)vpe_2_9(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[2][9]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[2][9]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[2][9]),
    .cast_data_o                                       (cast_data_pe_2_nw[2][9]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[2][9]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[2][9]),
    .merge_data_i                                      (merge_data_nw_2_pe[2][9]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[2][9]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[2][9]),
    .merge_data_o                                      (merge_data_pe_2_nw[2][9]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[2][9]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[2][9]),
    .gather_data_i                                     (gather_data_nw_2_pe[2][9]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[2][9]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[2][9]),
    .gather_data_o                                     (gather_data_pe_2_nw[2][9]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[2][9]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[2][9])
);


virtual_pe #(
    .cast_out                                          (cast_out_2_10),
    .merge_in                                          (merge_in_2_10),
    .merge_out                                         (merge_out_2_10),
    .gather_in                                         (gather_in_2_10),
    .gather_out                                        (gather_out_2_10),
    .x                                                 (2),
    .y                                                 (10)
)vpe_2_10(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[2][10]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[2][10]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[2][10]),
    .cast_data_o                                       (cast_data_pe_2_nw[2][10]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[2][10]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[2][10]),
    .merge_data_i                                      (merge_data_nw_2_pe[2][10]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[2][10]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[2][10]),
    .merge_data_o                                      (merge_data_pe_2_nw[2][10]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[2][10]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[2][10]),
    .gather_data_i                                     (gather_data_nw_2_pe[2][10]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[2][10]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[2][10]),
    .gather_data_o                                     (gather_data_pe_2_nw[2][10]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[2][10]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[2][10])
);


virtual_pe #(
    .cast_out                                          (cast_out_2_11),
    .merge_in                                          (merge_in_2_11),
    .merge_out                                         (merge_out_2_11),
    .gather_in                                         (gather_in_2_11),
    .gather_out                                        (gather_out_2_11),
    .x                                                 (2),
    .y                                                 (11)
)vpe_2_11(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[2][11]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[2][11]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[2][11]),
    .cast_data_o                                       (cast_data_pe_2_nw[2][11]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[2][11]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[2][11]),
    .merge_data_i                                      (merge_data_nw_2_pe[2][11]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[2][11]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[2][11]),
    .merge_data_o                                      (merge_data_pe_2_nw[2][11]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[2][11]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[2][11]),
    .gather_data_i                                     (gather_data_nw_2_pe[2][11]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[2][11]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[2][11]),
    .gather_data_o                                     (gather_data_pe_2_nw[2][11]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[2][11]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[2][11])
);


virtual_pe #(
    .cast_out                                          (cast_out_2_12),
    .merge_in                                          (merge_in_2_12),
    .merge_out                                         (merge_out_2_12),
    .gather_in                                         (gather_in_2_12),
    .gather_out                                        (gather_out_2_12),
    .x                                                 (2),
    .y                                                 (12)
)vpe_2_12(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[2][12]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[2][12]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[2][12]),
    .cast_data_o                                       (cast_data_pe_2_nw[2][12]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[2][12]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[2][12]),
    .merge_data_i                                      (merge_data_nw_2_pe[2][12]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[2][12]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[2][12]),
    .merge_data_o                                      (merge_data_pe_2_nw[2][12]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[2][12]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[2][12]),
    .gather_data_i                                     (gather_data_nw_2_pe[2][12]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[2][12]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[2][12]),
    .gather_data_o                                     (gather_data_pe_2_nw[2][12]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[2][12]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[2][12])
);


virtual_pe #(
    .cast_out                                          (cast_out_2_13),
    .merge_in                                          (merge_in_2_13),
    .merge_out                                         (merge_out_2_13),
    .gather_in                                         (gather_in_2_13),
    .gather_out                                        (gather_out_2_13),
    .x                                                 (2),
    .y                                                 (13)
)vpe_2_13(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[2][13]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[2][13]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[2][13]),
    .cast_data_o                                       (cast_data_pe_2_nw[2][13]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[2][13]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[2][13]),
    .merge_data_i                                      (merge_data_nw_2_pe[2][13]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[2][13]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[2][13]),
    .merge_data_o                                      (merge_data_pe_2_nw[2][13]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[2][13]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[2][13]),
    .gather_data_i                                     (gather_data_nw_2_pe[2][13]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[2][13]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[2][13]),
    .gather_data_o                                     (gather_data_pe_2_nw[2][13]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[2][13]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[2][13])
);


virtual_pe #(
    .cast_out                                          (cast_out_2_14),
    .merge_in                                          (merge_in_2_14),
    .merge_out                                         (merge_out_2_14),
    .gather_in                                         (gather_in_2_14),
    .gather_out                                        (gather_out_2_14),
    .x                                                 (2),
    .y                                                 (14)
)vpe_2_14(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[2][14]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[2][14]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[2][14]),
    .cast_data_o                                       (cast_data_pe_2_nw[2][14]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[2][14]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[2][14]),
    .merge_data_i                                      (merge_data_nw_2_pe[2][14]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[2][14]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[2][14]),
    .merge_data_o                                      (merge_data_pe_2_nw[2][14]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[2][14]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[2][14]),
    .gather_data_i                                     (gather_data_nw_2_pe[2][14]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[2][14]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[2][14]),
    .gather_data_o                                     (gather_data_pe_2_nw[2][14]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[2][14]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[2][14])
);


virtual_pe #(
    .cast_out                                          (cast_out_2_15),
    .merge_in                                          (merge_in_2_15),
    .merge_out                                         (merge_out_2_15),
    .gather_in                                         (gather_in_2_15),
    .gather_out                                        (gather_out_2_15),
    .x                                                 (2),
    .y                                                 (15)
)vpe_2_15(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[2][15]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[2][15]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[2][15]),
    .cast_data_o                                       (cast_data_pe_2_nw[2][15]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[2][15]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[2][15]),
    .merge_data_i                                      (merge_data_nw_2_pe[2][15]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[2][15]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[2][15]),
    .merge_data_o                                      (merge_data_pe_2_nw[2][15]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[2][15]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[2][15]),
    .gather_data_i                                     (gather_data_nw_2_pe[2][15]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[2][15]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[2][15]),
    .gather_data_o                                     (gather_data_pe_2_nw[2][15]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[2][15]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[2][15])
);


virtual_pe #(
    .cast_out                                          (cast_out_2_16),
    .merge_in                                          (merge_in_2_16),
    .merge_out                                         (merge_out_2_16),
    .gather_in                                         (gather_in_2_16),
    .gather_out                                        (gather_out_2_16),
    .x                                                 (2),
    .y                                                 (16)
)vpe_2_16(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[2][16]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[2][16]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[2][16]),
    .cast_data_o                                       (cast_data_pe_2_nw[2][16]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[2][16]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[2][16]),
    .merge_data_i                                      (merge_data_nw_2_pe[2][16]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[2][16]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[2][16]),
    .merge_data_o                                      (merge_data_pe_2_nw[2][16]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[2][16]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[2][16]),
    .gather_data_i                                     (gather_data_nw_2_pe[2][16]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[2][16]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[2][16]),
    .gather_data_o                                     (gather_data_pe_2_nw[2][16]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[2][16]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[2][16])
);


virtual_pe #(
    .cast_out                                          (cast_out_2_17),
    .merge_in                                          (merge_in_2_17),
    .merge_out                                         (merge_out_2_17),
    .gather_in                                         (gather_in_2_17),
    .gather_out                                        (gather_out_2_17),
    .x                                                 (2),
    .y                                                 (17)
)vpe_2_17(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[2][17]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[2][17]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[2][17]),
    .cast_data_o                                       (cast_data_pe_2_nw[2][17]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[2][17]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[2][17]),
    .merge_data_i                                      (merge_data_nw_2_pe[2][17]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[2][17]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[2][17]),
    .merge_data_o                                      (merge_data_pe_2_nw[2][17]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[2][17]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[2][17]),
    .gather_data_i                                     (gather_data_nw_2_pe[2][17]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[2][17]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[2][17]),
    .gather_data_o                                     (gather_data_pe_2_nw[2][17]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[2][17]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[2][17])
);


virtual_pe #(
    .cast_out                                          (cast_out_2_18),
    .merge_in                                          (merge_in_2_18),
    .merge_out                                         (merge_out_2_18),
    .gather_in                                         (gather_in_2_18),
    .gather_out                                        (gather_out_2_18),
    .x                                                 (2),
    .y                                                 (18)
)vpe_2_18(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[2][18]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[2][18]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[2][18]),
    .cast_data_o                                       (cast_data_pe_2_nw[2][18]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[2][18]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[2][18]),
    .merge_data_i                                      (merge_data_nw_2_pe[2][18]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[2][18]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[2][18]),
    .merge_data_o                                      (merge_data_pe_2_nw[2][18]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[2][18]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[2][18]),
    .gather_data_i                                     (gather_data_nw_2_pe[2][18]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[2][18]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[2][18]),
    .gather_data_o                                     (gather_data_pe_2_nw[2][18]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[2][18]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[2][18])
);


virtual_pe #(
    .cast_out                                          (cast_out_2_19),
    .merge_in                                          (merge_in_2_19),
    .merge_out                                         (merge_out_2_19),
    .gather_in                                         (gather_in_2_19),
    .gather_out                                        (gather_out_2_19),
    .x                                                 (2),
    .y                                                 (19)
)vpe_2_19(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[2][19]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[2][19]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[2][19]),
    .cast_data_o                                       (cast_data_pe_2_nw[2][19]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[2][19]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[2][19]),
    .merge_data_i                                      (merge_data_nw_2_pe[2][19]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[2][19]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[2][19]),
    .merge_data_o                                      (merge_data_pe_2_nw[2][19]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[2][19]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[2][19]),
    .gather_data_i                                     (gather_data_nw_2_pe[2][19]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[2][19]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[2][19]),
    .gather_data_o                                     (gather_data_pe_2_nw[2][19]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[2][19]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[2][19])
);


virtual_pe #(
    .cast_out                                          (cast_out_2_20),
    .merge_in                                          (merge_in_2_20),
    .merge_out                                         (merge_out_2_20),
    .gather_in                                         (gather_in_2_20),
    .gather_out                                        (gather_out_2_20),
    .x                                                 (2),
    .y                                                 (20)
)vpe_2_20(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[2][20]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[2][20]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[2][20]),
    .cast_data_o                                       (cast_data_pe_2_nw[2][20]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[2][20]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[2][20]),
    .merge_data_i                                      (merge_data_nw_2_pe[2][20]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[2][20]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[2][20]),
    .merge_data_o                                      (merge_data_pe_2_nw[2][20]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[2][20]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[2][20]),
    .gather_data_i                                     (gather_data_nw_2_pe[2][20]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[2][20]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[2][20]),
    .gather_data_o                                     (gather_data_pe_2_nw[2][20]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[2][20]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[2][20])
);


virtual_pe #(
    .cast_out                                          (cast_out_2_21),
    .merge_in                                          (merge_in_2_21),
    .merge_out                                         (merge_out_2_21),
    .gather_in                                         (gather_in_2_21),
    .gather_out                                        (gather_out_2_21),
    .x                                                 (2),
    .y                                                 (21)
)vpe_2_21(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[2][21]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[2][21]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[2][21]),
    .cast_data_o                                       (cast_data_pe_2_nw[2][21]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[2][21]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[2][21]),
    .merge_data_i                                      (merge_data_nw_2_pe[2][21]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[2][21]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[2][21]),
    .merge_data_o                                      (merge_data_pe_2_nw[2][21]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[2][21]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[2][21]),
    .gather_data_i                                     (gather_data_nw_2_pe[2][21]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[2][21]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[2][21]),
    .gather_data_o                                     (gather_data_pe_2_nw[2][21]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[2][21]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[2][21])
);


virtual_pe #(
    .cast_out                                          (cast_out_2_22),
    .merge_in                                          (merge_in_2_22),
    .merge_out                                         (merge_out_2_22),
    .gather_in                                         (gather_in_2_22),
    .gather_out                                        (gather_out_2_22),
    .x                                                 (2),
    .y                                                 (22)
)vpe_2_22(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[2][22]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[2][22]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[2][22]),
    .cast_data_o                                       (cast_data_pe_2_nw[2][22]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[2][22]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[2][22]),
    .merge_data_i                                      (merge_data_nw_2_pe[2][22]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[2][22]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[2][22]),
    .merge_data_o                                      (merge_data_pe_2_nw[2][22]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[2][22]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[2][22]),
    .gather_data_i                                     (gather_data_nw_2_pe[2][22]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[2][22]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[2][22]),
    .gather_data_o                                     (gather_data_pe_2_nw[2][22]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[2][22]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[2][22])
);


virtual_pe #(
    .cast_out                                          (cast_out_2_23),
    .merge_in                                          (merge_in_2_23),
    .merge_out                                         (merge_out_2_23),
    .gather_in                                         (gather_in_2_23),
    .gather_out                                        (gather_out_2_23),
    .x                                                 (2),
    .y                                                 (23)
)vpe_2_23(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[2][23]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[2][23]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[2][23]),
    .cast_data_o                                       (cast_data_pe_2_nw[2][23]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[2][23]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[2][23]),
    .merge_data_i                                      (merge_data_nw_2_pe[2][23]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[2][23]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[2][23]),
    .merge_data_o                                      (merge_data_pe_2_nw[2][23]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[2][23]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[2][23]),
    .gather_data_i                                     (gather_data_nw_2_pe[2][23]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[2][23]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[2][23]),
    .gather_data_o                                     (gather_data_pe_2_nw[2][23]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[2][23]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[2][23])
);


virtual_pe #(
    .cast_out                                          (cast_out_2_24),
    .merge_in                                          (merge_in_2_24),
    .merge_out                                         (merge_out_2_24),
    .gather_in                                         (gather_in_2_24),
    .gather_out                                        (gather_out_2_24),
    .x                                                 (2),
    .y                                                 (24)
)vpe_2_24(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[2][24]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[2][24]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[2][24]),
    .cast_data_o                                       (cast_data_pe_2_nw[2][24]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[2][24]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[2][24]),
    .merge_data_i                                      (merge_data_nw_2_pe[2][24]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[2][24]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[2][24]),
    .merge_data_o                                      (merge_data_pe_2_nw[2][24]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[2][24]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[2][24]),
    .gather_data_i                                     (gather_data_nw_2_pe[2][24]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[2][24]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[2][24]),
    .gather_data_o                                     (gather_data_pe_2_nw[2][24]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[2][24]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[2][24])
);


virtual_pe #(
    .cast_out                                          (cast_out_3_0),
    .merge_in                                          (merge_in_3_0),
    .merge_out                                         (merge_out_3_0),
    .gather_in                                         (gather_in_3_0),
    .gather_out                                        (gather_out_3_0),
    .x                                                 (3),
    .y                                                 (0)
)vpe_3_0(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[3][0]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[3][0]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[3][0]),
    .cast_data_o                                       (cast_data_pe_2_nw[3][0]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[3][0]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[3][0]),
    .merge_data_i                                      (merge_data_nw_2_pe[3][0]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[3][0]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[3][0]),
    .merge_data_o                                      (merge_data_pe_2_nw[3][0]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[3][0]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[3][0]),
    .gather_data_i                                     (gather_data_nw_2_pe[3][0]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[3][0]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[3][0]),
    .gather_data_o                                     (gather_data_pe_2_nw[3][0]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[3][0]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[3][0])
);


virtual_pe #(
    .cast_out                                          (cast_out_3_1),
    .merge_in                                          (merge_in_3_1),
    .merge_out                                         (merge_out_3_1),
    .gather_in                                         (gather_in_3_1),
    .gather_out                                        (gather_out_3_1),
    .x                                                 (3),
    .y                                                 (1)
)vpe_3_1(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[3][1]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[3][1]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[3][1]),
    .cast_data_o                                       (cast_data_pe_2_nw[3][1]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[3][1]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[3][1]),
    .merge_data_i                                      (merge_data_nw_2_pe[3][1]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[3][1]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[3][1]),
    .merge_data_o                                      (merge_data_pe_2_nw[3][1]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[3][1]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[3][1]),
    .gather_data_i                                     (gather_data_nw_2_pe[3][1]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[3][1]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[3][1]),
    .gather_data_o                                     (gather_data_pe_2_nw[3][1]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[3][1]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[3][1])
);


virtual_pe #(
    .cast_out                                          (cast_out_3_2),
    .merge_in                                          (merge_in_3_2),
    .merge_out                                         (merge_out_3_2),
    .gather_in                                         (gather_in_3_2),
    .gather_out                                        (gather_out_3_2),
    .x                                                 (3),
    .y                                                 (2)
)vpe_3_2(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[3][2]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[3][2]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[3][2]),
    .cast_data_o                                       (cast_data_pe_2_nw[3][2]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[3][2]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[3][2]),
    .merge_data_i                                      (merge_data_nw_2_pe[3][2]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[3][2]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[3][2]),
    .merge_data_o                                      (merge_data_pe_2_nw[3][2]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[3][2]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[3][2]),
    .gather_data_i                                     (gather_data_nw_2_pe[3][2]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[3][2]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[3][2]),
    .gather_data_o                                     (gather_data_pe_2_nw[3][2]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[3][2]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[3][2])
);


virtual_pe #(
    .cast_out                                          (cast_out_3_3),
    .merge_in                                          (merge_in_3_3),
    .merge_out                                         (merge_out_3_3),
    .gather_in                                         (gather_in_3_3),
    .gather_out                                        (gather_out_3_3),
    .x                                                 (3),
    .y                                                 (3)
)vpe_3_3(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[3][3]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[3][3]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[3][3]),
    .cast_data_o                                       (cast_data_pe_2_nw[3][3]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[3][3]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[3][3]),
    .merge_data_i                                      (merge_data_nw_2_pe[3][3]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[3][3]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[3][3]),
    .merge_data_o                                      (merge_data_pe_2_nw[3][3]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[3][3]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[3][3]),
    .gather_data_i                                     (gather_data_nw_2_pe[3][3]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[3][3]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[3][3]),
    .gather_data_o                                     (gather_data_pe_2_nw[3][3]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[3][3]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[3][3])
);


virtual_pe #(
    .cast_out                                          (cast_out_3_4),
    .merge_in                                          (merge_in_3_4),
    .merge_out                                         (merge_out_3_4),
    .gather_in                                         (gather_in_3_4),
    .gather_out                                        (gather_out_3_4),
    .x                                                 (3),
    .y                                                 (4)
)vpe_3_4(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[3][4]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[3][4]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[3][4]),
    .cast_data_o                                       (cast_data_pe_2_nw[3][4]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[3][4]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[3][4]),
    .merge_data_i                                      (merge_data_nw_2_pe[3][4]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[3][4]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[3][4]),
    .merge_data_o                                      (merge_data_pe_2_nw[3][4]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[3][4]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[3][4]),
    .gather_data_i                                     (gather_data_nw_2_pe[3][4]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[3][4]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[3][4]),
    .gather_data_o                                     (gather_data_pe_2_nw[3][4]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[3][4]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[3][4])
);


virtual_pe #(
    .cast_out                                          (cast_out_3_5),
    .merge_in                                          (merge_in_3_5),
    .merge_out                                         (merge_out_3_5),
    .gather_in                                         (gather_in_3_5),
    .gather_out                                        (gather_out_3_5),
    .x                                                 (3),
    .y                                                 (5)
)vpe_3_5(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[3][5]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[3][5]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[3][5]),
    .cast_data_o                                       (cast_data_pe_2_nw[3][5]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[3][5]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[3][5]),
    .merge_data_i                                      (merge_data_nw_2_pe[3][5]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[3][5]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[3][5]),
    .merge_data_o                                      (merge_data_pe_2_nw[3][5]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[3][5]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[3][5]),
    .gather_data_i                                     (gather_data_nw_2_pe[3][5]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[3][5]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[3][5]),
    .gather_data_o                                     (gather_data_pe_2_nw[3][5]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[3][5]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[3][5])
);


virtual_pe #(
    .cast_out                                          (cast_out_3_6),
    .merge_in                                          (merge_in_3_6),
    .merge_out                                         (merge_out_3_6),
    .gather_in                                         (gather_in_3_6),
    .gather_out                                        (gather_out_3_6),
    .x                                                 (3),
    .y                                                 (6)
)vpe_3_6(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[3][6]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[3][6]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[3][6]),
    .cast_data_o                                       (cast_data_pe_2_nw[3][6]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[3][6]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[3][6]),
    .merge_data_i                                      (merge_data_nw_2_pe[3][6]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[3][6]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[3][6]),
    .merge_data_o                                      (merge_data_pe_2_nw[3][6]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[3][6]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[3][6]),
    .gather_data_i                                     (gather_data_nw_2_pe[3][6]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[3][6]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[3][6]),
    .gather_data_o                                     (gather_data_pe_2_nw[3][6]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[3][6]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[3][6])
);


virtual_pe #(
    .cast_out                                          (cast_out_3_7),
    .merge_in                                          (merge_in_3_7),
    .merge_out                                         (merge_out_3_7),
    .gather_in                                         (gather_in_3_7),
    .gather_out                                        (gather_out_3_7),
    .x                                                 (3),
    .y                                                 (7)
)vpe_3_7(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[3][7]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[3][7]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[3][7]),
    .cast_data_o                                       (cast_data_pe_2_nw[3][7]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[3][7]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[3][7]),
    .merge_data_i                                      (merge_data_nw_2_pe[3][7]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[3][7]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[3][7]),
    .merge_data_o                                      (merge_data_pe_2_nw[3][7]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[3][7]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[3][7]),
    .gather_data_i                                     (gather_data_nw_2_pe[3][7]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[3][7]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[3][7]),
    .gather_data_o                                     (gather_data_pe_2_nw[3][7]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[3][7]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[3][7])
);


virtual_pe #(
    .cast_out                                          (cast_out_3_8),
    .merge_in                                          (merge_in_3_8),
    .merge_out                                         (merge_out_3_8),
    .gather_in                                         (gather_in_3_8),
    .gather_out                                        (gather_out_3_8),
    .x                                                 (3),
    .y                                                 (8)
)vpe_3_8(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[3][8]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[3][8]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[3][8]),
    .cast_data_o                                       (cast_data_pe_2_nw[3][8]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[3][8]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[3][8]),
    .merge_data_i                                      (merge_data_nw_2_pe[3][8]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[3][8]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[3][8]),
    .merge_data_o                                      (merge_data_pe_2_nw[3][8]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[3][8]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[3][8]),
    .gather_data_i                                     (gather_data_nw_2_pe[3][8]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[3][8]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[3][8]),
    .gather_data_o                                     (gather_data_pe_2_nw[3][8]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[3][8]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[3][8])
);


virtual_pe #(
    .cast_out                                          (cast_out_3_9),
    .merge_in                                          (merge_in_3_9),
    .merge_out                                         (merge_out_3_9),
    .gather_in                                         (gather_in_3_9),
    .gather_out                                        (gather_out_3_9),
    .x                                                 (3),
    .y                                                 (9)
)vpe_3_9(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[3][9]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[3][9]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[3][9]),
    .cast_data_o                                       (cast_data_pe_2_nw[3][9]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[3][9]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[3][9]),
    .merge_data_i                                      (merge_data_nw_2_pe[3][9]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[3][9]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[3][9]),
    .merge_data_o                                      (merge_data_pe_2_nw[3][9]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[3][9]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[3][9]),
    .gather_data_i                                     (gather_data_nw_2_pe[3][9]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[3][9]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[3][9]),
    .gather_data_o                                     (gather_data_pe_2_nw[3][9]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[3][9]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[3][9])
);


virtual_pe #(
    .cast_out                                          (cast_out_3_10),
    .merge_in                                          (merge_in_3_10),
    .merge_out                                         (merge_out_3_10),
    .gather_in                                         (gather_in_3_10),
    .gather_out                                        (gather_out_3_10),
    .x                                                 (3),
    .y                                                 (10)
)vpe_3_10(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[3][10]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[3][10]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[3][10]),
    .cast_data_o                                       (cast_data_pe_2_nw[3][10]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[3][10]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[3][10]),
    .merge_data_i                                      (merge_data_nw_2_pe[3][10]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[3][10]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[3][10]),
    .merge_data_o                                      (merge_data_pe_2_nw[3][10]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[3][10]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[3][10]),
    .gather_data_i                                     (gather_data_nw_2_pe[3][10]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[3][10]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[3][10]),
    .gather_data_o                                     (gather_data_pe_2_nw[3][10]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[3][10]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[3][10])
);


virtual_pe #(
    .cast_out                                          (cast_out_3_11),
    .merge_in                                          (merge_in_3_11),
    .merge_out                                         (merge_out_3_11),
    .gather_in                                         (gather_in_3_11),
    .gather_out                                        (gather_out_3_11),
    .x                                                 (3),
    .y                                                 (11)
)vpe_3_11(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[3][11]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[3][11]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[3][11]),
    .cast_data_o                                       (cast_data_pe_2_nw[3][11]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[3][11]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[3][11]),
    .merge_data_i                                      (merge_data_nw_2_pe[3][11]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[3][11]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[3][11]),
    .merge_data_o                                      (merge_data_pe_2_nw[3][11]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[3][11]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[3][11]),
    .gather_data_i                                     (gather_data_nw_2_pe[3][11]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[3][11]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[3][11]),
    .gather_data_o                                     (gather_data_pe_2_nw[3][11]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[3][11]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[3][11])
);


virtual_pe #(
    .cast_out                                          (cast_out_3_12),
    .merge_in                                          (merge_in_3_12),
    .merge_out                                         (merge_out_3_12),
    .gather_in                                         (gather_in_3_12),
    .gather_out                                        (gather_out_3_12),
    .x                                                 (3),
    .y                                                 (12)
)vpe_3_12(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[3][12]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[3][12]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[3][12]),
    .cast_data_o                                       (cast_data_pe_2_nw[3][12]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[3][12]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[3][12]),
    .merge_data_i                                      (merge_data_nw_2_pe[3][12]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[3][12]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[3][12]),
    .merge_data_o                                      (merge_data_pe_2_nw[3][12]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[3][12]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[3][12]),
    .gather_data_i                                     (gather_data_nw_2_pe[3][12]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[3][12]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[3][12]),
    .gather_data_o                                     (gather_data_pe_2_nw[3][12]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[3][12]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[3][12])
);


virtual_pe #(
    .cast_out                                          (cast_out_3_13),
    .merge_in                                          (merge_in_3_13),
    .merge_out                                         (merge_out_3_13),
    .gather_in                                         (gather_in_3_13),
    .gather_out                                        (gather_out_3_13),
    .x                                                 (3),
    .y                                                 (13)
)vpe_3_13(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[3][13]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[3][13]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[3][13]),
    .cast_data_o                                       (cast_data_pe_2_nw[3][13]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[3][13]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[3][13]),
    .merge_data_i                                      (merge_data_nw_2_pe[3][13]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[3][13]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[3][13]),
    .merge_data_o                                      (merge_data_pe_2_nw[3][13]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[3][13]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[3][13]),
    .gather_data_i                                     (gather_data_nw_2_pe[3][13]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[3][13]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[3][13]),
    .gather_data_o                                     (gather_data_pe_2_nw[3][13]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[3][13]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[3][13])
);


virtual_pe #(
    .cast_out                                          (cast_out_3_14),
    .merge_in                                          (merge_in_3_14),
    .merge_out                                         (merge_out_3_14),
    .gather_in                                         (gather_in_3_14),
    .gather_out                                        (gather_out_3_14),
    .x                                                 (3),
    .y                                                 (14)
)vpe_3_14(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[3][14]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[3][14]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[3][14]),
    .cast_data_o                                       (cast_data_pe_2_nw[3][14]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[3][14]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[3][14]),
    .merge_data_i                                      (merge_data_nw_2_pe[3][14]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[3][14]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[3][14]),
    .merge_data_o                                      (merge_data_pe_2_nw[3][14]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[3][14]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[3][14]),
    .gather_data_i                                     (gather_data_nw_2_pe[3][14]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[3][14]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[3][14]),
    .gather_data_o                                     (gather_data_pe_2_nw[3][14]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[3][14]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[3][14])
);


virtual_pe #(
    .cast_out                                          (cast_out_3_15),
    .merge_in                                          (merge_in_3_15),
    .merge_out                                         (merge_out_3_15),
    .gather_in                                         (gather_in_3_15),
    .gather_out                                        (gather_out_3_15),
    .x                                                 (3),
    .y                                                 (15)
)vpe_3_15(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[3][15]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[3][15]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[3][15]),
    .cast_data_o                                       (cast_data_pe_2_nw[3][15]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[3][15]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[3][15]),
    .merge_data_i                                      (merge_data_nw_2_pe[3][15]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[3][15]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[3][15]),
    .merge_data_o                                      (merge_data_pe_2_nw[3][15]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[3][15]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[3][15]),
    .gather_data_i                                     (gather_data_nw_2_pe[3][15]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[3][15]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[3][15]),
    .gather_data_o                                     (gather_data_pe_2_nw[3][15]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[3][15]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[3][15])
);


virtual_pe #(
    .cast_out                                          (cast_out_3_16),
    .merge_in                                          (merge_in_3_16),
    .merge_out                                         (merge_out_3_16),
    .gather_in                                         (gather_in_3_16),
    .gather_out                                        (gather_out_3_16),
    .x                                                 (3),
    .y                                                 (16)
)vpe_3_16(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[3][16]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[3][16]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[3][16]),
    .cast_data_o                                       (cast_data_pe_2_nw[3][16]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[3][16]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[3][16]),
    .merge_data_i                                      (merge_data_nw_2_pe[3][16]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[3][16]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[3][16]),
    .merge_data_o                                      (merge_data_pe_2_nw[3][16]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[3][16]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[3][16]),
    .gather_data_i                                     (gather_data_nw_2_pe[3][16]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[3][16]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[3][16]),
    .gather_data_o                                     (gather_data_pe_2_nw[3][16]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[3][16]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[3][16])
);


virtual_pe #(
    .cast_out                                          (cast_out_3_17),
    .merge_in                                          (merge_in_3_17),
    .merge_out                                         (merge_out_3_17),
    .gather_in                                         (gather_in_3_17),
    .gather_out                                        (gather_out_3_17),
    .x                                                 (3),
    .y                                                 (17)
)vpe_3_17(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[3][17]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[3][17]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[3][17]),
    .cast_data_o                                       (cast_data_pe_2_nw[3][17]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[3][17]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[3][17]),
    .merge_data_i                                      (merge_data_nw_2_pe[3][17]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[3][17]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[3][17]),
    .merge_data_o                                      (merge_data_pe_2_nw[3][17]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[3][17]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[3][17]),
    .gather_data_i                                     (gather_data_nw_2_pe[3][17]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[3][17]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[3][17]),
    .gather_data_o                                     (gather_data_pe_2_nw[3][17]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[3][17]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[3][17])
);


virtual_pe #(
    .cast_out                                          (cast_out_3_18),
    .merge_in                                          (merge_in_3_18),
    .merge_out                                         (merge_out_3_18),
    .gather_in                                         (gather_in_3_18),
    .gather_out                                        (gather_out_3_18),
    .x                                                 (3),
    .y                                                 (18)
)vpe_3_18(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[3][18]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[3][18]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[3][18]),
    .cast_data_o                                       (cast_data_pe_2_nw[3][18]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[3][18]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[3][18]),
    .merge_data_i                                      (merge_data_nw_2_pe[3][18]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[3][18]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[3][18]),
    .merge_data_o                                      (merge_data_pe_2_nw[3][18]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[3][18]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[3][18]),
    .gather_data_i                                     (gather_data_nw_2_pe[3][18]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[3][18]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[3][18]),
    .gather_data_o                                     (gather_data_pe_2_nw[3][18]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[3][18]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[3][18])
);


virtual_pe #(
    .cast_out                                          (cast_out_3_19),
    .merge_in                                          (merge_in_3_19),
    .merge_out                                         (merge_out_3_19),
    .gather_in                                         (gather_in_3_19),
    .gather_out                                        (gather_out_3_19),
    .x                                                 (3),
    .y                                                 (19)
)vpe_3_19(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[3][19]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[3][19]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[3][19]),
    .cast_data_o                                       (cast_data_pe_2_nw[3][19]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[3][19]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[3][19]),
    .merge_data_i                                      (merge_data_nw_2_pe[3][19]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[3][19]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[3][19]),
    .merge_data_o                                      (merge_data_pe_2_nw[3][19]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[3][19]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[3][19]),
    .gather_data_i                                     (gather_data_nw_2_pe[3][19]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[3][19]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[3][19]),
    .gather_data_o                                     (gather_data_pe_2_nw[3][19]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[3][19]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[3][19])
);


virtual_pe #(
    .cast_out                                          (cast_out_3_20),
    .merge_in                                          (merge_in_3_20),
    .merge_out                                         (merge_out_3_20),
    .gather_in                                         (gather_in_3_20),
    .gather_out                                        (gather_out_3_20),
    .x                                                 (3),
    .y                                                 (20)
)vpe_3_20(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[3][20]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[3][20]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[3][20]),
    .cast_data_o                                       (cast_data_pe_2_nw[3][20]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[3][20]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[3][20]),
    .merge_data_i                                      (merge_data_nw_2_pe[3][20]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[3][20]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[3][20]),
    .merge_data_o                                      (merge_data_pe_2_nw[3][20]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[3][20]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[3][20]),
    .gather_data_i                                     (gather_data_nw_2_pe[3][20]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[3][20]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[3][20]),
    .gather_data_o                                     (gather_data_pe_2_nw[3][20]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[3][20]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[3][20])
);


virtual_pe #(
    .cast_out                                          (cast_out_3_21),
    .merge_in                                          (merge_in_3_21),
    .merge_out                                         (merge_out_3_21),
    .gather_in                                         (gather_in_3_21),
    .gather_out                                        (gather_out_3_21),
    .x                                                 (3),
    .y                                                 (21)
)vpe_3_21(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[3][21]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[3][21]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[3][21]),
    .cast_data_o                                       (cast_data_pe_2_nw[3][21]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[3][21]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[3][21]),
    .merge_data_i                                      (merge_data_nw_2_pe[3][21]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[3][21]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[3][21]),
    .merge_data_o                                      (merge_data_pe_2_nw[3][21]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[3][21]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[3][21]),
    .gather_data_i                                     (gather_data_nw_2_pe[3][21]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[3][21]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[3][21]),
    .gather_data_o                                     (gather_data_pe_2_nw[3][21]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[3][21]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[3][21])
);


virtual_pe #(
    .cast_out                                          (cast_out_3_22),
    .merge_in                                          (merge_in_3_22),
    .merge_out                                         (merge_out_3_22),
    .gather_in                                         (gather_in_3_22),
    .gather_out                                        (gather_out_3_22),
    .x                                                 (3),
    .y                                                 (22)
)vpe_3_22(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[3][22]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[3][22]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[3][22]),
    .cast_data_o                                       (cast_data_pe_2_nw[3][22]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[3][22]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[3][22]),
    .merge_data_i                                      (merge_data_nw_2_pe[3][22]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[3][22]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[3][22]),
    .merge_data_o                                      (merge_data_pe_2_nw[3][22]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[3][22]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[3][22]),
    .gather_data_i                                     (gather_data_nw_2_pe[3][22]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[3][22]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[3][22]),
    .gather_data_o                                     (gather_data_pe_2_nw[3][22]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[3][22]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[3][22])
);


virtual_pe #(
    .cast_out                                          (cast_out_3_23),
    .merge_in                                          (merge_in_3_23),
    .merge_out                                         (merge_out_3_23),
    .gather_in                                         (gather_in_3_23),
    .gather_out                                        (gather_out_3_23),
    .x                                                 (3),
    .y                                                 (23)
)vpe_3_23(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[3][23]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[3][23]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[3][23]),
    .cast_data_o                                       (cast_data_pe_2_nw[3][23]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[3][23]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[3][23]),
    .merge_data_i                                      (merge_data_nw_2_pe[3][23]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[3][23]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[3][23]),
    .merge_data_o                                      (merge_data_pe_2_nw[3][23]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[3][23]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[3][23]),
    .gather_data_i                                     (gather_data_nw_2_pe[3][23]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[3][23]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[3][23]),
    .gather_data_o                                     (gather_data_pe_2_nw[3][23]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[3][23]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[3][23])
);


virtual_pe #(
    .cast_out                                          (cast_out_3_24),
    .merge_in                                          (merge_in_3_24),
    .merge_out                                         (merge_out_3_24),
    .gather_in                                         (gather_in_3_24),
    .gather_out                                        (gather_out_3_24),
    .x                                                 (3),
    .y                                                 (24)
)vpe_3_24(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[3][24]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[3][24]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[3][24]),
    .cast_data_o                                       (cast_data_pe_2_nw[3][24]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[3][24]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[3][24]),
    .merge_data_i                                      (merge_data_nw_2_pe[3][24]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[3][24]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[3][24]),
    .merge_data_o                                      (merge_data_pe_2_nw[3][24]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[3][24]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[3][24]),
    .gather_data_i                                     (gather_data_nw_2_pe[3][24]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[3][24]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[3][24]),
    .gather_data_o                                     (gather_data_pe_2_nw[3][24]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[3][24]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[3][24])
);


virtual_pe #(
    .cast_out                                          (cast_out_4_0),
    .merge_in                                          (merge_in_4_0),
    .merge_out                                         (merge_out_4_0),
    .gather_in                                         (gather_in_4_0),
    .gather_out                                        (gather_out_4_0),
    .x                                                 (4),
    .y                                                 (0)
)vpe_4_0(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[4][0]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[4][0]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[4][0]),
    .cast_data_o                                       (cast_data_pe_2_nw[4][0]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[4][0]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[4][0]),
    .merge_data_i                                      (merge_data_nw_2_pe[4][0]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[4][0]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[4][0]),
    .merge_data_o                                      (merge_data_pe_2_nw[4][0]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[4][0]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[4][0]),
    .gather_data_i                                     (gather_data_nw_2_pe[4][0]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[4][0]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[4][0]),
    .gather_data_o                                     (gather_data_pe_2_nw[4][0]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[4][0]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[4][0])
);


virtual_pe #(
    .cast_out                                          (cast_out_4_1),
    .merge_in                                          (merge_in_4_1),
    .merge_out                                         (merge_out_4_1),
    .gather_in                                         (gather_in_4_1),
    .gather_out                                        (gather_out_4_1),
    .x                                                 (4),
    .y                                                 (1)
)vpe_4_1(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[4][1]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[4][1]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[4][1]),
    .cast_data_o                                       (cast_data_pe_2_nw[4][1]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[4][1]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[4][1]),
    .merge_data_i                                      (merge_data_nw_2_pe[4][1]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[4][1]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[4][1]),
    .merge_data_o                                      (merge_data_pe_2_nw[4][1]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[4][1]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[4][1]),
    .gather_data_i                                     (gather_data_nw_2_pe[4][1]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[4][1]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[4][1]),
    .gather_data_o                                     (gather_data_pe_2_nw[4][1]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[4][1]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[4][1])
);


virtual_pe #(
    .cast_out                                          (cast_out_4_2),
    .merge_in                                          (merge_in_4_2),
    .merge_out                                         (merge_out_4_2),
    .gather_in                                         (gather_in_4_2),
    .gather_out                                        (gather_out_4_2),
    .x                                                 (4),
    .y                                                 (2)
)vpe_4_2(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[4][2]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[4][2]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[4][2]),
    .cast_data_o                                       (cast_data_pe_2_nw[4][2]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[4][2]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[4][2]),
    .merge_data_i                                      (merge_data_nw_2_pe[4][2]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[4][2]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[4][2]),
    .merge_data_o                                      (merge_data_pe_2_nw[4][2]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[4][2]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[4][2]),
    .gather_data_i                                     (gather_data_nw_2_pe[4][2]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[4][2]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[4][2]),
    .gather_data_o                                     (gather_data_pe_2_nw[4][2]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[4][2]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[4][2])
);


virtual_pe #(
    .cast_out                                          (cast_out_4_3),
    .merge_in                                          (merge_in_4_3),
    .merge_out                                         (merge_out_4_3),
    .gather_in                                         (gather_in_4_3),
    .gather_out                                        (gather_out_4_3),
    .x                                                 (4),
    .y                                                 (3)
)vpe_4_3(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[4][3]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[4][3]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[4][3]),
    .cast_data_o                                       (cast_data_pe_2_nw[4][3]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[4][3]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[4][3]),
    .merge_data_i                                      (merge_data_nw_2_pe[4][3]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[4][3]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[4][3]),
    .merge_data_o                                      (merge_data_pe_2_nw[4][3]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[4][3]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[4][3]),
    .gather_data_i                                     (gather_data_nw_2_pe[4][3]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[4][3]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[4][3]),
    .gather_data_o                                     (gather_data_pe_2_nw[4][3]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[4][3]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[4][3])
);


virtual_pe #(
    .cast_out                                          (cast_out_4_4),
    .merge_in                                          (merge_in_4_4),
    .merge_out                                         (merge_out_4_4),
    .gather_in                                         (gather_in_4_4),
    .gather_out                                        (gather_out_4_4),
    .x                                                 (4),
    .y                                                 (4)
)vpe_4_4(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[4][4]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[4][4]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[4][4]),
    .cast_data_o                                       (cast_data_pe_2_nw[4][4]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[4][4]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[4][4]),
    .merge_data_i                                      (merge_data_nw_2_pe[4][4]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[4][4]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[4][4]),
    .merge_data_o                                      (merge_data_pe_2_nw[4][4]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[4][4]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[4][4]),
    .gather_data_i                                     (gather_data_nw_2_pe[4][4]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[4][4]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[4][4]),
    .gather_data_o                                     (gather_data_pe_2_nw[4][4]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[4][4]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[4][4])
);


virtual_pe #(
    .cast_out                                          (cast_out_4_5),
    .merge_in                                          (merge_in_4_5),
    .merge_out                                         (merge_out_4_5),
    .gather_in                                         (gather_in_4_5),
    .gather_out                                        (gather_out_4_5),
    .x                                                 (4),
    .y                                                 (5)
)vpe_4_5(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[4][5]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[4][5]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[4][5]),
    .cast_data_o                                       (cast_data_pe_2_nw[4][5]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[4][5]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[4][5]),
    .merge_data_i                                      (merge_data_nw_2_pe[4][5]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[4][5]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[4][5]),
    .merge_data_o                                      (merge_data_pe_2_nw[4][5]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[4][5]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[4][5]),
    .gather_data_i                                     (gather_data_nw_2_pe[4][5]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[4][5]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[4][5]),
    .gather_data_o                                     (gather_data_pe_2_nw[4][5]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[4][5]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[4][5])
);


virtual_pe #(
    .cast_out                                          (cast_out_4_6),
    .merge_in                                          (merge_in_4_6),
    .merge_out                                         (merge_out_4_6),
    .gather_in                                         (gather_in_4_6),
    .gather_out                                        (gather_out_4_6),
    .x                                                 (4),
    .y                                                 (6)
)vpe_4_6(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[4][6]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[4][6]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[4][6]),
    .cast_data_o                                       (cast_data_pe_2_nw[4][6]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[4][6]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[4][6]),
    .merge_data_i                                      (merge_data_nw_2_pe[4][6]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[4][6]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[4][6]),
    .merge_data_o                                      (merge_data_pe_2_nw[4][6]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[4][6]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[4][6]),
    .gather_data_i                                     (gather_data_nw_2_pe[4][6]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[4][6]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[4][6]),
    .gather_data_o                                     (gather_data_pe_2_nw[4][6]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[4][6]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[4][6])
);


virtual_pe #(
    .cast_out                                          (cast_out_4_7),
    .merge_in                                          (merge_in_4_7),
    .merge_out                                         (merge_out_4_7),
    .gather_in                                         (gather_in_4_7),
    .gather_out                                        (gather_out_4_7),
    .x                                                 (4),
    .y                                                 (7)
)vpe_4_7(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[4][7]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[4][7]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[4][7]),
    .cast_data_o                                       (cast_data_pe_2_nw[4][7]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[4][7]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[4][7]),
    .merge_data_i                                      (merge_data_nw_2_pe[4][7]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[4][7]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[4][7]),
    .merge_data_o                                      (merge_data_pe_2_nw[4][7]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[4][7]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[4][7]),
    .gather_data_i                                     (gather_data_nw_2_pe[4][7]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[4][7]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[4][7]),
    .gather_data_o                                     (gather_data_pe_2_nw[4][7]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[4][7]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[4][7])
);


virtual_pe #(
    .cast_out                                          (cast_out_4_8),
    .merge_in                                          (merge_in_4_8),
    .merge_out                                         (merge_out_4_8),
    .gather_in                                         (gather_in_4_8),
    .gather_out                                        (gather_out_4_8),
    .x                                                 (4),
    .y                                                 (8)
)vpe_4_8(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[4][8]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[4][8]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[4][8]),
    .cast_data_o                                       (cast_data_pe_2_nw[4][8]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[4][8]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[4][8]),
    .merge_data_i                                      (merge_data_nw_2_pe[4][8]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[4][8]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[4][8]),
    .merge_data_o                                      (merge_data_pe_2_nw[4][8]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[4][8]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[4][8]),
    .gather_data_i                                     (gather_data_nw_2_pe[4][8]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[4][8]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[4][8]),
    .gather_data_o                                     (gather_data_pe_2_nw[4][8]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[4][8]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[4][8])
);


virtual_pe #(
    .cast_out                                          (cast_out_4_9),
    .merge_in                                          (merge_in_4_9),
    .merge_out                                         (merge_out_4_9),
    .gather_in                                         (gather_in_4_9),
    .gather_out                                        (gather_out_4_9),
    .x                                                 (4),
    .y                                                 (9)
)vpe_4_9(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[4][9]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[4][9]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[4][9]),
    .cast_data_o                                       (cast_data_pe_2_nw[4][9]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[4][9]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[4][9]),
    .merge_data_i                                      (merge_data_nw_2_pe[4][9]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[4][9]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[4][9]),
    .merge_data_o                                      (merge_data_pe_2_nw[4][9]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[4][9]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[4][9]),
    .gather_data_i                                     (gather_data_nw_2_pe[4][9]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[4][9]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[4][9]),
    .gather_data_o                                     (gather_data_pe_2_nw[4][9]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[4][9]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[4][9])
);


virtual_pe #(
    .cast_out                                          (cast_out_4_10),
    .merge_in                                          (merge_in_4_10),
    .merge_out                                         (merge_out_4_10),
    .gather_in                                         (gather_in_4_10),
    .gather_out                                        (gather_out_4_10),
    .x                                                 (4),
    .y                                                 (10)
)vpe_4_10(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[4][10]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[4][10]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[4][10]),
    .cast_data_o                                       (cast_data_pe_2_nw[4][10]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[4][10]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[4][10]),
    .merge_data_i                                      (merge_data_nw_2_pe[4][10]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[4][10]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[4][10]),
    .merge_data_o                                      (merge_data_pe_2_nw[4][10]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[4][10]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[4][10]),
    .gather_data_i                                     (gather_data_nw_2_pe[4][10]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[4][10]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[4][10]),
    .gather_data_o                                     (gather_data_pe_2_nw[4][10]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[4][10]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[4][10])
);


virtual_pe #(
    .cast_out                                          (cast_out_4_11),
    .merge_in                                          (merge_in_4_11),
    .merge_out                                         (merge_out_4_11),
    .gather_in                                         (gather_in_4_11),
    .gather_out                                        (gather_out_4_11),
    .x                                                 (4),
    .y                                                 (11)
)vpe_4_11(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[4][11]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[4][11]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[4][11]),
    .cast_data_o                                       (cast_data_pe_2_nw[4][11]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[4][11]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[4][11]),
    .merge_data_i                                      (merge_data_nw_2_pe[4][11]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[4][11]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[4][11]),
    .merge_data_o                                      (merge_data_pe_2_nw[4][11]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[4][11]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[4][11]),
    .gather_data_i                                     (gather_data_nw_2_pe[4][11]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[4][11]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[4][11]),
    .gather_data_o                                     (gather_data_pe_2_nw[4][11]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[4][11]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[4][11])
);


virtual_pe #(
    .cast_out                                          (cast_out_4_12),
    .merge_in                                          (merge_in_4_12),
    .merge_out                                         (merge_out_4_12),
    .gather_in                                         (gather_in_4_12),
    .gather_out                                        (gather_out_4_12),
    .x                                                 (4),
    .y                                                 (12)
)vpe_4_12(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[4][12]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[4][12]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[4][12]),
    .cast_data_o                                       (cast_data_pe_2_nw[4][12]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[4][12]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[4][12]),
    .merge_data_i                                      (merge_data_nw_2_pe[4][12]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[4][12]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[4][12]),
    .merge_data_o                                      (merge_data_pe_2_nw[4][12]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[4][12]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[4][12]),
    .gather_data_i                                     (gather_data_nw_2_pe[4][12]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[4][12]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[4][12]),
    .gather_data_o                                     (gather_data_pe_2_nw[4][12]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[4][12]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[4][12])
);


virtual_pe #(
    .cast_out                                          (cast_out_4_13),
    .merge_in                                          (merge_in_4_13),
    .merge_out                                         (merge_out_4_13),
    .gather_in                                         (gather_in_4_13),
    .gather_out                                        (gather_out_4_13),
    .x                                                 (4),
    .y                                                 (13)
)vpe_4_13(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[4][13]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[4][13]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[4][13]),
    .cast_data_o                                       (cast_data_pe_2_nw[4][13]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[4][13]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[4][13]),
    .merge_data_i                                      (merge_data_nw_2_pe[4][13]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[4][13]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[4][13]),
    .merge_data_o                                      (merge_data_pe_2_nw[4][13]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[4][13]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[4][13]),
    .gather_data_i                                     (gather_data_nw_2_pe[4][13]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[4][13]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[4][13]),
    .gather_data_o                                     (gather_data_pe_2_nw[4][13]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[4][13]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[4][13])
);


virtual_pe #(
    .cast_out                                          (cast_out_4_14),
    .merge_in                                          (merge_in_4_14),
    .merge_out                                         (merge_out_4_14),
    .gather_in                                         (gather_in_4_14),
    .gather_out                                        (gather_out_4_14),
    .x                                                 (4),
    .y                                                 (14)
)vpe_4_14(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[4][14]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[4][14]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[4][14]),
    .cast_data_o                                       (cast_data_pe_2_nw[4][14]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[4][14]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[4][14]),
    .merge_data_i                                      (merge_data_nw_2_pe[4][14]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[4][14]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[4][14]),
    .merge_data_o                                      (merge_data_pe_2_nw[4][14]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[4][14]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[4][14]),
    .gather_data_i                                     (gather_data_nw_2_pe[4][14]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[4][14]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[4][14]),
    .gather_data_o                                     (gather_data_pe_2_nw[4][14]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[4][14]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[4][14])
);


virtual_pe #(
    .cast_out                                          (cast_out_4_15),
    .merge_in                                          (merge_in_4_15),
    .merge_out                                         (merge_out_4_15),
    .gather_in                                         (gather_in_4_15),
    .gather_out                                        (gather_out_4_15),
    .x                                                 (4),
    .y                                                 (15)
)vpe_4_15(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[4][15]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[4][15]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[4][15]),
    .cast_data_o                                       (cast_data_pe_2_nw[4][15]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[4][15]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[4][15]),
    .merge_data_i                                      (merge_data_nw_2_pe[4][15]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[4][15]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[4][15]),
    .merge_data_o                                      (merge_data_pe_2_nw[4][15]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[4][15]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[4][15]),
    .gather_data_i                                     (gather_data_nw_2_pe[4][15]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[4][15]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[4][15]),
    .gather_data_o                                     (gather_data_pe_2_nw[4][15]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[4][15]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[4][15])
);


virtual_pe #(
    .cast_out                                          (cast_out_4_16),
    .merge_in                                          (merge_in_4_16),
    .merge_out                                         (merge_out_4_16),
    .gather_in                                         (gather_in_4_16),
    .gather_out                                        (gather_out_4_16),
    .x                                                 (4),
    .y                                                 (16)
)vpe_4_16(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[4][16]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[4][16]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[4][16]),
    .cast_data_o                                       (cast_data_pe_2_nw[4][16]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[4][16]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[4][16]),
    .merge_data_i                                      (merge_data_nw_2_pe[4][16]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[4][16]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[4][16]),
    .merge_data_o                                      (merge_data_pe_2_nw[4][16]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[4][16]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[4][16]),
    .gather_data_i                                     (gather_data_nw_2_pe[4][16]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[4][16]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[4][16]),
    .gather_data_o                                     (gather_data_pe_2_nw[4][16]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[4][16]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[4][16])
);


virtual_pe #(
    .cast_out                                          (cast_out_4_17),
    .merge_in                                          (merge_in_4_17),
    .merge_out                                         (merge_out_4_17),
    .gather_in                                         (gather_in_4_17),
    .gather_out                                        (gather_out_4_17),
    .x                                                 (4),
    .y                                                 (17)
)vpe_4_17(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[4][17]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[4][17]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[4][17]),
    .cast_data_o                                       (cast_data_pe_2_nw[4][17]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[4][17]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[4][17]),
    .merge_data_i                                      (merge_data_nw_2_pe[4][17]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[4][17]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[4][17]),
    .merge_data_o                                      (merge_data_pe_2_nw[4][17]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[4][17]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[4][17]),
    .gather_data_i                                     (gather_data_nw_2_pe[4][17]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[4][17]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[4][17]),
    .gather_data_o                                     (gather_data_pe_2_nw[4][17]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[4][17]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[4][17])
);


virtual_pe #(
    .cast_out                                          (cast_out_4_18),
    .merge_in                                          (merge_in_4_18),
    .merge_out                                         (merge_out_4_18),
    .gather_in                                         (gather_in_4_18),
    .gather_out                                        (gather_out_4_18),
    .x                                                 (4),
    .y                                                 (18)
)vpe_4_18(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[4][18]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[4][18]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[4][18]),
    .cast_data_o                                       (cast_data_pe_2_nw[4][18]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[4][18]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[4][18]),
    .merge_data_i                                      (merge_data_nw_2_pe[4][18]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[4][18]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[4][18]),
    .merge_data_o                                      (merge_data_pe_2_nw[4][18]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[4][18]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[4][18]),
    .gather_data_i                                     (gather_data_nw_2_pe[4][18]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[4][18]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[4][18]),
    .gather_data_o                                     (gather_data_pe_2_nw[4][18]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[4][18]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[4][18])
);


virtual_pe #(
    .cast_out                                          (cast_out_4_19),
    .merge_in                                          (merge_in_4_19),
    .merge_out                                         (merge_out_4_19),
    .gather_in                                         (gather_in_4_19),
    .gather_out                                        (gather_out_4_19),
    .x                                                 (4),
    .y                                                 (19)
)vpe_4_19(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[4][19]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[4][19]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[4][19]),
    .cast_data_o                                       (cast_data_pe_2_nw[4][19]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[4][19]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[4][19]),
    .merge_data_i                                      (merge_data_nw_2_pe[4][19]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[4][19]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[4][19]),
    .merge_data_o                                      (merge_data_pe_2_nw[4][19]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[4][19]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[4][19]),
    .gather_data_i                                     (gather_data_nw_2_pe[4][19]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[4][19]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[4][19]),
    .gather_data_o                                     (gather_data_pe_2_nw[4][19]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[4][19]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[4][19])
);


virtual_pe #(
    .cast_out                                          (cast_out_4_20),
    .merge_in                                          (merge_in_4_20),
    .merge_out                                         (merge_out_4_20),
    .gather_in                                         (gather_in_4_20),
    .gather_out                                        (gather_out_4_20),
    .x                                                 (4),
    .y                                                 (20)
)vpe_4_20(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[4][20]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[4][20]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[4][20]),
    .cast_data_o                                       (cast_data_pe_2_nw[4][20]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[4][20]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[4][20]),
    .merge_data_i                                      (merge_data_nw_2_pe[4][20]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[4][20]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[4][20]),
    .merge_data_o                                      (merge_data_pe_2_nw[4][20]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[4][20]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[4][20]),
    .gather_data_i                                     (gather_data_nw_2_pe[4][20]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[4][20]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[4][20]),
    .gather_data_o                                     (gather_data_pe_2_nw[4][20]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[4][20]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[4][20])
);


virtual_pe #(
    .cast_out                                          (cast_out_4_21),
    .merge_in                                          (merge_in_4_21),
    .merge_out                                         (merge_out_4_21),
    .gather_in                                         (gather_in_4_21),
    .gather_out                                        (gather_out_4_21),
    .x                                                 (4),
    .y                                                 (21)
)vpe_4_21(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[4][21]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[4][21]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[4][21]),
    .cast_data_o                                       (cast_data_pe_2_nw[4][21]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[4][21]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[4][21]),
    .merge_data_i                                      (merge_data_nw_2_pe[4][21]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[4][21]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[4][21]),
    .merge_data_o                                      (merge_data_pe_2_nw[4][21]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[4][21]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[4][21]),
    .gather_data_i                                     (gather_data_nw_2_pe[4][21]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[4][21]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[4][21]),
    .gather_data_o                                     (gather_data_pe_2_nw[4][21]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[4][21]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[4][21])
);


virtual_pe #(
    .cast_out                                          (cast_out_4_22),
    .merge_in                                          (merge_in_4_22),
    .merge_out                                         (merge_out_4_22),
    .gather_in                                         (gather_in_4_22),
    .gather_out                                        (gather_out_4_22),
    .x                                                 (4),
    .y                                                 (22)
)vpe_4_22(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[4][22]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[4][22]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[4][22]),
    .cast_data_o                                       (cast_data_pe_2_nw[4][22]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[4][22]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[4][22]),
    .merge_data_i                                      (merge_data_nw_2_pe[4][22]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[4][22]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[4][22]),
    .merge_data_o                                      (merge_data_pe_2_nw[4][22]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[4][22]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[4][22]),
    .gather_data_i                                     (gather_data_nw_2_pe[4][22]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[4][22]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[4][22]),
    .gather_data_o                                     (gather_data_pe_2_nw[4][22]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[4][22]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[4][22])
);


virtual_pe #(
    .cast_out                                          (cast_out_4_23),
    .merge_in                                          (merge_in_4_23),
    .merge_out                                         (merge_out_4_23),
    .gather_in                                         (gather_in_4_23),
    .gather_out                                        (gather_out_4_23),
    .x                                                 (4),
    .y                                                 (23)
)vpe_4_23(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[4][23]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[4][23]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[4][23]),
    .cast_data_o                                       (cast_data_pe_2_nw[4][23]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[4][23]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[4][23]),
    .merge_data_i                                      (merge_data_nw_2_pe[4][23]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[4][23]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[4][23]),
    .merge_data_o                                      (merge_data_pe_2_nw[4][23]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[4][23]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[4][23]),
    .gather_data_i                                     (gather_data_nw_2_pe[4][23]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[4][23]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[4][23]),
    .gather_data_o                                     (gather_data_pe_2_nw[4][23]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[4][23]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[4][23])
);


virtual_pe #(
    .cast_out                                          (cast_out_4_24),
    .merge_in                                          (merge_in_4_24),
    .merge_out                                         (merge_out_4_24),
    .gather_in                                         (gather_in_4_24),
    .gather_out                                        (gather_out_4_24),
    .x                                                 (4),
    .y                                                 (24)
)vpe_4_24(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[4][24]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[4][24]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[4][24]),
    .cast_data_o                                       (cast_data_pe_2_nw[4][24]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[4][24]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[4][24]),
    .merge_data_i                                      (merge_data_nw_2_pe[4][24]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[4][24]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[4][24]),
    .merge_data_o                                      (merge_data_pe_2_nw[4][24]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[4][24]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[4][24]),
    .gather_data_i                                     (gather_data_nw_2_pe[4][24]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[4][24]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[4][24]),
    .gather_data_o                                     (gather_data_pe_2_nw[4][24]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[4][24]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[4][24])
);


virtual_pe #(
    .cast_out                                          (cast_out_5_0),
    .merge_in                                          (merge_in_5_0),
    .merge_out                                         (merge_out_5_0),
    .gather_in                                         (gather_in_5_0),
    .gather_out                                        (gather_out_5_0),
    .x                                                 (5),
    .y                                                 (0)
)vpe_5_0(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[5][0]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[5][0]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[5][0]),
    .cast_data_o                                       (cast_data_pe_2_nw[5][0]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[5][0]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[5][0]),
    .merge_data_i                                      (merge_data_nw_2_pe[5][0]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[5][0]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[5][0]),
    .merge_data_o                                      (merge_data_pe_2_nw[5][0]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[5][0]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[5][0]),
    .gather_data_i                                     (gather_data_nw_2_pe[5][0]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[5][0]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[5][0]),
    .gather_data_o                                     (gather_data_pe_2_nw[5][0]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[5][0]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[5][0])
);


virtual_pe #(
    .cast_out                                          (cast_out_5_1),
    .merge_in                                          (merge_in_5_1),
    .merge_out                                         (merge_out_5_1),
    .gather_in                                         (gather_in_5_1),
    .gather_out                                        (gather_out_5_1),
    .x                                                 (5),
    .y                                                 (1)
)vpe_5_1(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[5][1]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[5][1]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[5][1]),
    .cast_data_o                                       (cast_data_pe_2_nw[5][1]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[5][1]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[5][1]),
    .merge_data_i                                      (merge_data_nw_2_pe[5][1]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[5][1]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[5][1]),
    .merge_data_o                                      (merge_data_pe_2_nw[5][1]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[5][1]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[5][1]),
    .gather_data_i                                     (gather_data_nw_2_pe[5][1]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[5][1]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[5][1]),
    .gather_data_o                                     (gather_data_pe_2_nw[5][1]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[5][1]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[5][1])
);


virtual_pe #(
    .cast_out                                          (cast_out_5_2),
    .merge_in                                          (merge_in_5_2),
    .merge_out                                         (merge_out_5_2),
    .gather_in                                         (gather_in_5_2),
    .gather_out                                        (gather_out_5_2),
    .x                                                 (5),
    .y                                                 (2)
)vpe_5_2(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[5][2]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[5][2]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[5][2]),
    .cast_data_o                                       (cast_data_pe_2_nw[5][2]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[5][2]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[5][2]),
    .merge_data_i                                      (merge_data_nw_2_pe[5][2]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[5][2]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[5][2]),
    .merge_data_o                                      (merge_data_pe_2_nw[5][2]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[5][2]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[5][2]),
    .gather_data_i                                     (gather_data_nw_2_pe[5][2]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[5][2]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[5][2]),
    .gather_data_o                                     (gather_data_pe_2_nw[5][2]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[5][2]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[5][2])
);


virtual_pe #(
    .cast_out                                          (cast_out_5_3),
    .merge_in                                          (merge_in_5_3),
    .merge_out                                         (merge_out_5_3),
    .gather_in                                         (gather_in_5_3),
    .gather_out                                        (gather_out_5_3),
    .x                                                 (5),
    .y                                                 (3)
)vpe_5_3(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[5][3]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[5][3]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[5][3]),
    .cast_data_o                                       (cast_data_pe_2_nw[5][3]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[5][3]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[5][3]),
    .merge_data_i                                      (merge_data_nw_2_pe[5][3]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[5][3]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[5][3]),
    .merge_data_o                                      (merge_data_pe_2_nw[5][3]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[5][3]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[5][3]),
    .gather_data_i                                     (gather_data_nw_2_pe[5][3]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[5][3]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[5][3]),
    .gather_data_o                                     (gather_data_pe_2_nw[5][3]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[5][3]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[5][3])
);


virtual_pe #(
    .cast_out                                          (cast_out_5_4),
    .merge_in                                          (merge_in_5_4),
    .merge_out                                         (merge_out_5_4),
    .gather_in                                         (gather_in_5_4),
    .gather_out                                        (gather_out_5_4),
    .x                                                 (5),
    .y                                                 (4)
)vpe_5_4(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[5][4]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[5][4]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[5][4]),
    .cast_data_o                                       (cast_data_pe_2_nw[5][4]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[5][4]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[5][4]),
    .merge_data_i                                      (merge_data_nw_2_pe[5][4]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[5][4]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[5][4]),
    .merge_data_o                                      (merge_data_pe_2_nw[5][4]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[5][4]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[5][4]),
    .gather_data_i                                     (gather_data_nw_2_pe[5][4]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[5][4]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[5][4]),
    .gather_data_o                                     (gather_data_pe_2_nw[5][4]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[5][4]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[5][4])
);


virtual_pe #(
    .cast_out                                          (cast_out_5_5),
    .merge_in                                          (merge_in_5_5),
    .merge_out                                         (merge_out_5_5),
    .gather_in                                         (gather_in_5_5),
    .gather_out                                        (gather_out_5_5),
    .x                                                 (5),
    .y                                                 (5)
)vpe_5_5(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[5][5]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[5][5]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[5][5]),
    .cast_data_o                                       (cast_data_pe_2_nw[5][5]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[5][5]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[5][5]),
    .merge_data_i                                      (merge_data_nw_2_pe[5][5]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[5][5]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[5][5]),
    .merge_data_o                                      (merge_data_pe_2_nw[5][5]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[5][5]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[5][5]),
    .gather_data_i                                     (gather_data_nw_2_pe[5][5]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[5][5]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[5][5]),
    .gather_data_o                                     (gather_data_pe_2_nw[5][5]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[5][5]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[5][5])
);


virtual_pe #(
    .cast_out                                          (cast_out_5_6),
    .merge_in                                          (merge_in_5_6),
    .merge_out                                         (merge_out_5_6),
    .gather_in                                         (gather_in_5_6),
    .gather_out                                        (gather_out_5_6),
    .x                                                 (5),
    .y                                                 (6)
)vpe_5_6(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[5][6]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[5][6]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[5][6]),
    .cast_data_o                                       (cast_data_pe_2_nw[5][6]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[5][6]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[5][6]),
    .merge_data_i                                      (merge_data_nw_2_pe[5][6]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[5][6]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[5][6]),
    .merge_data_o                                      (merge_data_pe_2_nw[5][6]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[5][6]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[5][6]),
    .gather_data_i                                     (gather_data_nw_2_pe[5][6]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[5][6]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[5][6]),
    .gather_data_o                                     (gather_data_pe_2_nw[5][6]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[5][6]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[5][6])
);


virtual_pe #(
    .cast_out                                          (cast_out_5_7),
    .merge_in                                          (merge_in_5_7),
    .merge_out                                         (merge_out_5_7),
    .gather_in                                         (gather_in_5_7),
    .gather_out                                        (gather_out_5_7),
    .x                                                 (5),
    .y                                                 (7)
)vpe_5_7(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[5][7]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[5][7]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[5][7]),
    .cast_data_o                                       (cast_data_pe_2_nw[5][7]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[5][7]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[5][7]),
    .merge_data_i                                      (merge_data_nw_2_pe[5][7]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[5][7]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[5][7]),
    .merge_data_o                                      (merge_data_pe_2_nw[5][7]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[5][7]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[5][7]),
    .gather_data_i                                     (gather_data_nw_2_pe[5][7]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[5][7]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[5][7]),
    .gather_data_o                                     (gather_data_pe_2_nw[5][7]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[5][7]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[5][7])
);


virtual_pe #(
    .cast_out                                          (cast_out_5_8),
    .merge_in                                          (merge_in_5_8),
    .merge_out                                         (merge_out_5_8),
    .gather_in                                         (gather_in_5_8),
    .gather_out                                        (gather_out_5_8),
    .x                                                 (5),
    .y                                                 (8)
)vpe_5_8(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[5][8]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[5][8]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[5][8]),
    .cast_data_o                                       (cast_data_pe_2_nw[5][8]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[5][8]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[5][8]),
    .merge_data_i                                      (merge_data_nw_2_pe[5][8]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[5][8]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[5][8]),
    .merge_data_o                                      (merge_data_pe_2_nw[5][8]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[5][8]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[5][8]),
    .gather_data_i                                     (gather_data_nw_2_pe[5][8]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[5][8]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[5][8]),
    .gather_data_o                                     (gather_data_pe_2_nw[5][8]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[5][8]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[5][8])
);


virtual_pe #(
    .cast_out                                          (cast_out_5_9),
    .merge_in                                          (merge_in_5_9),
    .merge_out                                         (merge_out_5_9),
    .gather_in                                         (gather_in_5_9),
    .gather_out                                        (gather_out_5_9),
    .x                                                 (5),
    .y                                                 (9)
)vpe_5_9(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[5][9]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[5][9]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[5][9]),
    .cast_data_o                                       (cast_data_pe_2_nw[5][9]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[5][9]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[5][9]),
    .merge_data_i                                      (merge_data_nw_2_pe[5][9]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[5][9]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[5][9]),
    .merge_data_o                                      (merge_data_pe_2_nw[5][9]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[5][9]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[5][9]),
    .gather_data_i                                     (gather_data_nw_2_pe[5][9]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[5][9]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[5][9]),
    .gather_data_o                                     (gather_data_pe_2_nw[5][9]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[5][9]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[5][9])
);


virtual_pe #(
    .cast_out                                          (cast_out_5_10),
    .merge_in                                          (merge_in_5_10),
    .merge_out                                         (merge_out_5_10),
    .gather_in                                         (gather_in_5_10),
    .gather_out                                        (gather_out_5_10),
    .x                                                 (5),
    .y                                                 (10)
)vpe_5_10(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[5][10]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[5][10]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[5][10]),
    .cast_data_o                                       (cast_data_pe_2_nw[5][10]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[5][10]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[5][10]),
    .merge_data_i                                      (merge_data_nw_2_pe[5][10]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[5][10]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[5][10]),
    .merge_data_o                                      (merge_data_pe_2_nw[5][10]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[5][10]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[5][10]),
    .gather_data_i                                     (gather_data_nw_2_pe[5][10]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[5][10]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[5][10]),
    .gather_data_o                                     (gather_data_pe_2_nw[5][10]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[5][10]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[5][10])
);


virtual_pe #(
    .cast_out                                          (cast_out_5_11),
    .merge_in                                          (merge_in_5_11),
    .merge_out                                         (merge_out_5_11),
    .gather_in                                         (gather_in_5_11),
    .gather_out                                        (gather_out_5_11),
    .x                                                 (5),
    .y                                                 (11)
)vpe_5_11(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[5][11]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[5][11]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[5][11]),
    .cast_data_o                                       (cast_data_pe_2_nw[5][11]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[5][11]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[5][11]),
    .merge_data_i                                      (merge_data_nw_2_pe[5][11]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[5][11]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[5][11]),
    .merge_data_o                                      (merge_data_pe_2_nw[5][11]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[5][11]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[5][11]),
    .gather_data_i                                     (gather_data_nw_2_pe[5][11]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[5][11]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[5][11]),
    .gather_data_o                                     (gather_data_pe_2_nw[5][11]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[5][11]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[5][11])
);


virtual_pe #(
    .cast_out                                          (cast_out_5_12),
    .merge_in                                          (merge_in_5_12),
    .merge_out                                         (merge_out_5_12),
    .gather_in                                         (gather_in_5_12),
    .gather_out                                        (gather_out_5_12),
    .x                                                 (5),
    .y                                                 (12)
)vpe_5_12(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[5][12]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[5][12]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[5][12]),
    .cast_data_o                                       (cast_data_pe_2_nw[5][12]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[5][12]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[5][12]),
    .merge_data_i                                      (merge_data_nw_2_pe[5][12]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[5][12]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[5][12]),
    .merge_data_o                                      (merge_data_pe_2_nw[5][12]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[5][12]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[5][12]),
    .gather_data_i                                     (gather_data_nw_2_pe[5][12]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[5][12]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[5][12]),
    .gather_data_o                                     (gather_data_pe_2_nw[5][12]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[5][12]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[5][12])
);


virtual_pe #(
    .cast_out                                          (cast_out_5_13),
    .merge_in                                          (merge_in_5_13),
    .merge_out                                         (merge_out_5_13),
    .gather_in                                         (gather_in_5_13),
    .gather_out                                        (gather_out_5_13),
    .x                                                 (5),
    .y                                                 (13)
)vpe_5_13(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[5][13]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[5][13]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[5][13]),
    .cast_data_o                                       (cast_data_pe_2_nw[5][13]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[5][13]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[5][13]),
    .merge_data_i                                      (merge_data_nw_2_pe[5][13]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[5][13]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[5][13]),
    .merge_data_o                                      (merge_data_pe_2_nw[5][13]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[5][13]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[5][13]),
    .gather_data_i                                     (gather_data_nw_2_pe[5][13]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[5][13]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[5][13]),
    .gather_data_o                                     (gather_data_pe_2_nw[5][13]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[5][13]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[5][13])
);


virtual_pe #(
    .cast_out                                          (cast_out_5_14),
    .merge_in                                          (merge_in_5_14),
    .merge_out                                         (merge_out_5_14),
    .gather_in                                         (gather_in_5_14),
    .gather_out                                        (gather_out_5_14),
    .x                                                 (5),
    .y                                                 (14)
)vpe_5_14(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[5][14]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[5][14]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[5][14]),
    .cast_data_o                                       (cast_data_pe_2_nw[5][14]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[5][14]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[5][14]),
    .merge_data_i                                      (merge_data_nw_2_pe[5][14]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[5][14]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[5][14]),
    .merge_data_o                                      (merge_data_pe_2_nw[5][14]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[5][14]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[5][14]),
    .gather_data_i                                     (gather_data_nw_2_pe[5][14]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[5][14]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[5][14]),
    .gather_data_o                                     (gather_data_pe_2_nw[5][14]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[5][14]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[5][14])
);


virtual_pe #(
    .cast_out                                          (cast_out_5_15),
    .merge_in                                          (merge_in_5_15),
    .merge_out                                         (merge_out_5_15),
    .gather_in                                         (gather_in_5_15),
    .gather_out                                        (gather_out_5_15),
    .x                                                 (5),
    .y                                                 (15)
)vpe_5_15(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[5][15]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[5][15]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[5][15]),
    .cast_data_o                                       (cast_data_pe_2_nw[5][15]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[5][15]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[5][15]),
    .merge_data_i                                      (merge_data_nw_2_pe[5][15]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[5][15]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[5][15]),
    .merge_data_o                                      (merge_data_pe_2_nw[5][15]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[5][15]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[5][15]),
    .gather_data_i                                     (gather_data_nw_2_pe[5][15]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[5][15]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[5][15]),
    .gather_data_o                                     (gather_data_pe_2_nw[5][15]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[5][15]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[5][15])
);


virtual_pe #(
    .cast_out                                          (cast_out_5_16),
    .merge_in                                          (merge_in_5_16),
    .merge_out                                         (merge_out_5_16),
    .gather_in                                         (gather_in_5_16),
    .gather_out                                        (gather_out_5_16),
    .x                                                 (5),
    .y                                                 (16)
)vpe_5_16(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[5][16]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[5][16]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[5][16]),
    .cast_data_o                                       (cast_data_pe_2_nw[5][16]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[5][16]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[5][16]),
    .merge_data_i                                      (merge_data_nw_2_pe[5][16]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[5][16]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[5][16]),
    .merge_data_o                                      (merge_data_pe_2_nw[5][16]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[5][16]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[5][16]),
    .gather_data_i                                     (gather_data_nw_2_pe[5][16]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[5][16]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[5][16]),
    .gather_data_o                                     (gather_data_pe_2_nw[5][16]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[5][16]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[5][16])
);


virtual_pe #(
    .cast_out                                          (cast_out_5_17),
    .merge_in                                          (merge_in_5_17),
    .merge_out                                         (merge_out_5_17),
    .gather_in                                         (gather_in_5_17),
    .gather_out                                        (gather_out_5_17),
    .x                                                 (5),
    .y                                                 (17)
)vpe_5_17(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[5][17]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[5][17]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[5][17]),
    .cast_data_o                                       (cast_data_pe_2_nw[5][17]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[5][17]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[5][17]),
    .merge_data_i                                      (merge_data_nw_2_pe[5][17]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[5][17]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[5][17]),
    .merge_data_o                                      (merge_data_pe_2_nw[5][17]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[5][17]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[5][17]),
    .gather_data_i                                     (gather_data_nw_2_pe[5][17]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[5][17]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[5][17]),
    .gather_data_o                                     (gather_data_pe_2_nw[5][17]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[5][17]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[5][17])
);


virtual_pe #(
    .cast_out                                          (cast_out_5_18),
    .merge_in                                          (merge_in_5_18),
    .merge_out                                         (merge_out_5_18),
    .gather_in                                         (gather_in_5_18),
    .gather_out                                        (gather_out_5_18),
    .x                                                 (5),
    .y                                                 (18)
)vpe_5_18(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[5][18]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[5][18]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[5][18]),
    .cast_data_o                                       (cast_data_pe_2_nw[5][18]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[5][18]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[5][18]),
    .merge_data_i                                      (merge_data_nw_2_pe[5][18]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[5][18]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[5][18]),
    .merge_data_o                                      (merge_data_pe_2_nw[5][18]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[5][18]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[5][18]),
    .gather_data_i                                     (gather_data_nw_2_pe[5][18]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[5][18]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[5][18]),
    .gather_data_o                                     (gather_data_pe_2_nw[5][18]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[5][18]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[5][18])
);


virtual_pe #(
    .cast_out                                          (cast_out_5_19),
    .merge_in                                          (merge_in_5_19),
    .merge_out                                         (merge_out_5_19),
    .gather_in                                         (gather_in_5_19),
    .gather_out                                        (gather_out_5_19),
    .x                                                 (5),
    .y                                                 (19)
)vpe_5_19(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[5][19]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[5][19]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[5][19]),
    .cast_data_o                                       (cast_data_pe_2_nw[5][19]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[5][19]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[5][19]),
    .merge_data_i                                      (merge_data_nw_2_pe[5][19]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[5][19]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[5][19]),
    .merge_data_o                                      (merge_data_pe_2_nw[5][19]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[5][19]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[5][19]),
    .gather_data_i                                     (gather_data_nw_2_pe[5][19]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[5][19]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[5][19]),
    .gather_data_o                                     (gather_data_pe_2_nw[5][19]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[5][19]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[5][19])
);


virtual_pe #(
    .cast_out                                          (cast_out_5_20),
    .merge_in                                          (merge_in_5_20),
    .merge_out                                         (merge_out_5_20),
    .gather_in                                         (gather_in_5_20),
    .gather_out                                        (gather_out_5_20),
    .x                                                 (5),
    .y                                                 (20)
)vpe_5_20(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[5][20]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[5][20]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[5][20]),
    .cast_data_o                                       (cast_data_pe_2_nw[5][20]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[5][20]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[5][20]),
    .merge_data_i                                      (merge_data_nw_2_pe[5][20]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[5][20]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[5][20]),
    .merge_data_o                                      (merge_data_pe_2_nw[5][20]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[5][20]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[5][20]),
    .gather_data_i                                     (gather_data_nw_2_pe[5][20]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[5][20]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[5][20]),
    .gather_data_o                                     (gather_data_pe_2_nw[5][20]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[5][20]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[5][20])
);


virtual_pe #(
    .cast_out                                          (cast_out_5_21),
    .merge_in                                          (merge_in_5_21),
    .merge_out                                         (merge_out_5_21),
    .gather_in                                         (gather_in_5_21),
    .gather_out                                        (gather_out_5_21),
    .x                                                 (5),
    .y                                                 (21)
)vpe_5_21(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[5][21]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[5][21]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[5][21]),
    .cast_data_o                                       (cast_data_pe_2_nw[5][21]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[5][21]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[5][21]),
    .merge_data_i                                      (merge_data_nw_2_pe[5][21]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[5][21]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[5][21]),
    .merge_data_o                                      (merge_data_pe_2_nw[5][21]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[5][21]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[5][21]),
    .gather_data_i                                     (gather_data_nw_2_pe[5][21]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[5][21]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[5][21]),
    .gather_data_o                                     (gather_data_pe_2_nw[5][21]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[5][21]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[5][21])
);


virtual_pe #(
    .cast_out                                          (cast_out_5_22),
    .merge_in                                          (merge_in_5_22),
    .merge_out                                         (merge_out_5_22),
    .gather_in                                         (gather_in_5_22),
    .gather_out                                        (gather_out_5_22),
    .x                                                 (5),
    .y                                                 (22)
)vpe_5_22(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[5][22]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[5][22]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[5][22]),
    .cast_data_o                                       (cast_data_pe_2_nw[5][22]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[5][22]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[5][22]),
    .merge_data_i                                      (merge_data_nw_2_pe[5][22]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[5][22]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[5][22]),
    .merge_data_o                                      (merge_data_pe_2_nw[5][22]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[5][22]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[5][22]),
    .gather_data_i                                     (gather_data_nw_2_pe[5][22]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[5][22]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[5][22]),
    .gather_data_o                                     (gather_data_pe_2_nw[5][22]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[5][22]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[5][22])
);


virtual_pe #(
    .cast_out                                          (cast_out_5_23),
    .merge_in                                          (merge_in_5_23),
    .merge_out                                         (merge_out_5_23),
    .gather_in                                         (gather_in_5_23),
    .gather_out                                        (gather_out_5_23),
    .x                                                 (5),
    .y                                                 (23)
)vpe_5_23(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[5][23]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[5][23]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[5][23]),
    .cast_data_o                                       (cast_data_pe_2_nw[5][23]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[5][23]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[5][23]),
    .merge_data_i                                      (merge_data_nw_2_pe[5][23]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[5][23]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[5][23]),
    .merge_data_o                                      (merge_data_pe_2_nw[5][23]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[5][23]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[5][23]),
    .gather_data_i                                     (gather_data_nw_2_pe[5][23]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[5][23]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[5][23]),
    .gather_data_o                                     (gather_data_pe_2_nw[5][23]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[5][23]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[5][23])
);


virtual_pe #(
    .cast_out                                          (cast_out_5_24),
    .merge_in                                          (merge_in_5_24),
    .merge_out                                         (merge_out_5_24),
    .gather_in                                         (gather_in_5_24),
    .gather_out                                        (gather_out_5_24),
    .x                                                 (5),
    .y                                                 (24)
)vpe_5_24(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[5][24]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[5][24]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[5][24]),
    .cast_data_o                                       (cast_data_pe_2_nw[5][24]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[5][24]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[5][24]),
    .merge_data_i                                      (merge_data_nw_2_pe[5][24]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[5][24]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[5][24]),
    .merge_data_o                                      (merge_data_pe_2_nw[5][24]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[5][24]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[5][24]),
    .gather_data_i                                     (gather_data_nw_2_pe[5][24]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[5][24]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[5][24]),
    .gather_data_o                                     (gather_data_pe_2_nw[5][24]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[5][24]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[5][24])
);


virtual_pe #(
    .cast_out                                          (cast_out_6_0),
    .merge_in                                          (merge_in_6_0),
    .merge_out                                         (merge_out_6_0),
    .gather_in                                         (gather_in_6_0),
    .gather_out                                        (gather_out_6_0),
    .x                                                 (6),
    .y                                                 (0)
)vpe_6_0(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[6][0]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[6][0]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[6][0]),
    .cast_data_o                                       (cast_data_pe_2_nw[6][0]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[6][0]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[6][0]),
    .merge_data_i                                      (merge_data_nw_2_pe[6][0]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[6][0]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[6][0]),
    .merge_data_o                                      (merge_data_pe_2_nw[6][0]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[6][0]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[6][0]),
    .gather_data_i                                     (gather_data_nw_2_pe[6][0]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[6][0]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[6][0]),
    .gather_data_o                                     (gather_data_pe_2_nw[6][0]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[6][0]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[6][0])
);


virtual_pe #(
    .cast_out                                          (cast_out_6_1),
    .merge_in                                          (merge_in_6_1),
    .merge_out                                         (merge_out_6_1),
    .gather_in                                         (gather_in_6_1),
    .gather_out                                        (gather_out_6_1),
    .x                                                 (6),
    .y                                                 (1)
)vpe_6_1(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[6][1]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[6][1]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[6][1]),
    .cast_data_o                                       (cast_data_pe_2_nw[6][1]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[6][1]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[6][1]),
    .merge_data_i                                      (merge_data_nw_2_pe[6][1]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[6][1]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[6][1]),
    .merge_data_o                                      (merge_data_pe_2_nw[6][1]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[6][1]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[6][1]),
    .gather_data_i                                     (gather_data_nw_2_pe[6][1]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[6][1]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[6][1]),
    .gather_data_o                                     (gather_data_pe_2_nw[6][1]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[6][1]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[6][1])
);


virtual_pe #(
    .cast_out                                          (cast_out_6_2),
    .merge_in                                          (merge_in_6_2),
    .merge_out                                         (merge_out_6_2),
    .gather_in                                         (gather_in_6_2),
    .gather_out                                        (gather_out_6_2),
    .x                                                 (6),
    .y                                                 (2)
)vpe_6_2(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[6][2]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[6][2]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[6][2]),
    .cast_data_o                                       (cast_data_pe_2_nw[6][2]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[6][2]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[6][2]),
    .merge_data_i                                      (merge_data_nw_2_pe[6][2]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[6][2]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[6][2]),
    .merge_data_o                                      (merge_data_pe_2_nw[6][2]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[6][2]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[6][2]),
    .gather_data_i                                     (gather_data_nw_2_pe[6][2]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[6][2]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[6][2]),
    .gather_data_o                                     (gather_data_pe_2_nw[6][2]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[6][2]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[6][2])
);


virtual_pe #(
    .cast_out                                          (cast_out_6_3),
    .merge_in                                          (merge_in_6_3),
    .merge_out                                         (merge_out_6_3),
    .gather_in                                         (gather_in_6_3),
    .gather_out                                        (gather_out_6_3),
    .x                                                 (6),
    .y                                                 (3)
)vpe_6_3(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[6][3]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[6][3]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[6][3]),
    .cast_data_o                                       (cast_data_pe_2_nw[6][3]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[6][3]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[6][3]),
    .merge_data_i                                      (merge_data_nw_2_pe[6][3]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[6][3]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[6][3]),
    .merge_data_o                                      (merge_data_pe_2_nw[6][3]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[6][3]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[6][3]),
    .gather_data_i                                     (gather_data_nw_2_pe[6][3]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[6][3]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[6][3]),
    .gather_data_o                                     (gather_data_pe_2_nw[6][3]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[6][3]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[6][3])
);


virtual_pe #(
    .cast_out                                          (cast_out_6_4),
    .merge_in                                          (merge_in_6_4),
    .merge_out                                         (merge_out_6_4),
    .gather_in                                         (gather_in_6_4),
    .gather_out                                        (gather_out_6_4),
    .x                                                 (6),
    .y                                                 (4)
)vpe_6_4(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[6][4]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[6][4]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[6][4]),
    .cast_data_o                                       (cast_data_pe_2_nw[6][4]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[6][4]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[6][4]),
    .merge_data_i                                      (merge_data_nw_2_pe[6][4]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[6][4]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[6][4]),
    .merge_data_o                                      (merge_data_pe_2_nw[6][4]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[6][4]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[6][4]),
    .gather_data_i                                     (gather_data_nw_2_pe[6][4]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[6][4]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[6][4]),
    .gather_data_o                                     (gather_data_pe_2_nw[6][4]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[6][4]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[6][4])
);


virtual_pe #(
    .cast_out                                          (cast_out_6_5),
    .merge_in                                          (merge_in_6_5),
    .merge_out                                         (merge_out_6_5),
    .gather_in                                         (gather_in_6_5),
    .gather_out                                        (gather_out_6_5),
    .x                                                 (6),
    .y                                                 (5)
)vpe_6_5(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[6][5]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[6][5]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[6][5]),
    .cast_data_o                                       (cast_data_pe_2_nw[6][5]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[6][5]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[6][5]),
    .merge_data_i                                      (merge_data_nw_2_pe[6][5]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[6][5]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[6][5]),
    .merge_data_o                                      (merge_data_pe_2_nw[6][5]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[6][5]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[6][5]),
    .gather_data_i                                     (gather_data_nw_2_pe[6][5]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[6][5]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[6][5]),
    .gather_data_o                                     (gather_data_pe_2_nw[6][5]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[6][5]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[6][5])
);


virtual_pe #(
    .cast_out                                          (cast_out_6_6),
    .merge_in                                          (merge_in_6_6),
    .merge_out                                         (merge_out_6_6),
    .gather_in                                         (gather_in_6_6),
    .gather_out                                        (gather_out_6_6),
    .x                                                 (6),
    .y                                                 (6)
)vpe_6_6(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[6][6]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[6][6]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[6][6]),
    .cast_data_o                                       (cast_data_pe_2_nw[6][6]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[6][6]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[6][6]),
    .merge_data_i                                      (merge_data_nw_2_pe[6][6]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[6][6]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[6][6]),
    .merge_data_o                                      (merge_data_pe_2_nw[6][6]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[6][6]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[6][6]),
    .gather_data_i                                     (gather_data_nw_2_pe[6][6]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[6][6]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[6][6]),
    .gather_data_o                                     (gather_data_pe_2_nw[6][6]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[6][6]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[6][6])
);


virtual_pe #(
    .cast_out                                          (cast_out_6_7),
    .merge_in                                          (merge_in_6_7),
    .merge_out                                         (merge_out_6_7),
    .gather_in                                         (gather_in_6_7),
    .gather_out                                        (gather_out_6_7),
    .x                                                 (6),
    .y                                                 (7)
)vpe_6_7(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[6][7]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[6][7]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[6][7]),
    .cast_data_o                                       (cast_data_pe_2_nw[6][7]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[6][7]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[6][7]),
    .merge_data_i                                      (merge_data_nw_2_pe[6][7]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[6][7]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[6][7]),
    .merge_data_o                                      (merge_data_pe_2_nw[6][7]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[6][7]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[6][7]),
    .gather_data_i                                     (gather_data_nw_2_pe[6][7]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[6][7]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[6][7]),
    .gather_data_o                                     (gather_data_pe_2_nw[6][7]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[6][7]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[6][7])
);


virtual_pe #(
    .cast_out                                          (cast_out_6_8),
    .merge_in                                          (merge_in_6_8),
    .merge_out                                         (merge_out_6_8),
    .gather_in                                         (gather_in_6_8),
    .gather_out                                        (gather_out_6_8),
    .x                                                 (6),
    .y                                                 (8)
)vpe_6_8(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[6][8]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[6][8]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[6][8]),
    .cast_data_o                                       (cast_data_pe_2_nw[6][8]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[6][8]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[6][8]),
    .merge_data_i                                      (merge_data_nw_2_pe[6][8]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[6][8]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[6][8]),
    .merge_data_o                                      (merge_data_pe_2_nw[6][8]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[6][8]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[6][8]),
    .gather_data_i                                     (gather_data_nw_2_pe[6][8]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[6][8]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[6][8]),
    .gather_data_o                                     (gather_data_pe_2_nw[6][8]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[6][8]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[6][8])
);


virtual_pe #(
    .cast_out                                          (cast_out_6_9),
    .merge_in                                          (merge_in_6_9),
    .merge_out                                         (merge_out_6_9),
    .gather_in                                         (gather_in_6_9),
    .gather_out                                        (gather_out_6_9),
    .x                                                 (6),
    .y                                                 (9)
)vpe_6_9(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[6][9]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[6][9]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[6][9]),
    .cast_data_o                                       (cast_data_pe_2_nw[6][9]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[6][9]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[6][9]),
    .merge_data_i                                      (merge_data_nw_2_pe[6][9]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[6][9]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[6][9]),
    .merge_data_o                                      (merge_data_pe_2_nw[6][9]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[6][9]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[6][9]),
    .gather_data_i                                     (gather_data_nw_2_pe[6][9]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[6][9]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[6][9]),
    .gather_data_o                                     (gather_data_pe_2_nw[6][9]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[6][9]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[6][9])
);


virtual_pe #(
    .cast_out                                          (cast_out_6_10),
    .merge_in                                          (merge_in_6_10),
    .merge_out                                         (merge_out_6_10),
    .gather_in                                         (gather_in_6_10),
    .gather_out                                        (gather_out_6_10),
    .x                                                 (6),
    .y                                                 (10)
)vpe_6_10(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[6][10]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[6][10]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[6][10]),
    .cast_data_o                                       (cast_data_pe_2_nw[6][10]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[6][10]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[6][10]),
    .merge_data_i                                      (merge_data_nw_2_pe[6][10]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[6][10]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[6][10]),
    .merge_data_o                                      (merge_data_pe_2_nw[6][10]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[6][10]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[6][10]),
    .gather_data_i                                     (gather_data_nw_2_pe[6][10]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[6][10]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[6][10]),
    .gather_data_o                                     (gather_data_pe_2_nw[6][10]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[6][10]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[6][10])
);


virtual_pe #(
    .cast_out                                          (cast_out_6_11),
    .merge_in                                          (merge_in_6_11),
    .merge_out                                         (merge_out_6_11),
    .gather_in                                         (gather_in_6_11),
    .gather_out                                        (gather_out_6_11),
    .x                                                 (6),
    .y                                                 (11)
)vpe_6_11(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[6][11]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[6][11]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[6][11]),
    .cast_data_o                                       (cast_data_pe_2_nw[6][11]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[6][11]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[6][11]),
    .merge_data_i                                      (merge_data_nw_2_pe[6][11]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[6][11]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[6][11]),
    .merge_data_o                                      (merge_data_pe_2_nw[6][11]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[6][11]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[6][11]),
    .gather_data_i                                     (gather_data_nw_2_pe[6][11]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[6][11]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[6][11]),
    .gather_data_o                                     (gather_data_pe_2_nw[6][11]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[6][11]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[6][11])
);


virtual_pe #(
    .cast_out                                          (cast_out_6_12),
    .merge_in                                          (merge_in_6_12),
    .merge_out                                         (merge_out_6_12),
    .gather_in                                         (gather_in_6_12),
    .gather_out                                        (gather_out_6_12),
    .x                                                 (6),
    .y                                                 (12)
)vpe_6_12(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[6][12]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[6][12]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[6][12]),
    .cast_data_o                                       (cast_data_pe_2_nw[6][12]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[6][12]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[6][12]),
    .merge_data_i                                      (merge_data_nw_2_pe[6][12]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[6][12]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[6][12]),
    .merge_data_o                                      (merge_data_pe_2_nw[6][12]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[6][12]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[6][12]),
    .gather_data_i                                     (gather_data_nw_2_pe[6][12]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[6][12]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[6][12]),
    .gather_data_o                                     (gather_data_pe_2_nw[6][12]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[6][12]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[6][12])
);


virtual_pe #(
    .cast_out                                          (cast_out_6_13),
    .merge_in                                          (merge_in_6_13),
    .merge_out                                         (merge_out_6_13),
    .gather_in                                         (gather_in_6_13),
    .gather_out                                        (gather_out_6_13),
    .x                                                 (6),
    .y                                                 (13)
)vpe_6_13(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[6][13]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[6][13]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[6][13]),
    .cast_data_o                                       (cast_data_pe_2_nw[6][13]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[6][13]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[6][13]),
    .merge_data_i                                      (merge_data_nw_2_pe[6][13]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[6][13]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[6][13]),
    .merge_data_o                                      (merge_data_pe_2_nw[6][13]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[6][13]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[6][13]),
    .gather_data_i                                     (gather_data_nw_2_pe[6][13]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[6][13]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[6][13]),
    .gather_data_o                                     (gather_data_pe_2_nw[6][13]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[6][13]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[6][13])
);


virtual_pe #(
    .cast_out                                          (cast_out_6_14),
    .merge_in                                          (merge_in_6_14),
    .merge_out                                         (merge_out_6_14),
    .gather_in                                         (gather_in_6_14),
    .gather_out                                        (gather_out_6_14),
    .x                                                 (6),
    .y                                                 (14)
)vpe_6_14(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[6][14]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[6][14]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[6][14]),
    .cast_data_o                                       (cast_data_pe_2_nw[6][14]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[6][14]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[6][14]),
    .merge_data_i                                      (merge_data_nw_2_pe[6][14]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[6][14]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[6][14]),
    .merge_data_o                                      (merge_data_pe_2_nw[6][14]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[6][14]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[6][14]),
    .gather_data_i                                     (gather_data_nw_2_pe[6][14]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[6][14]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[6][14]),
    .gather_data_o                                     (gather_data_pe_2_nw[6][14]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[6][14]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[6][14])
);


virtual_pe #(
    .cast_out                                          (cast_out_6_15),
    .merge_in                                          (merge_in_6_15),
    .merge_out                                         (merge_out_6_15),
    .gather_in                                         (gather_in_6_15),
    .gather_out                                        (gather_out_6_15),
    .x                                                 (6),
    .y                                                 (15)
)vpe_6_15(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[6][15]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[6][15]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[6][15]),
    .cast_data_o                                       (cast_data_pe_2_nw[6][15]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[6][15]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[6][15]),
    .merge_data_i                                      (merge_data_nw_2_pe[6][15]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[6][15]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[6][15]),
    .merge_data_o                                      (merge_data_pe_2_nw[6][15]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[6][15]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[6][15]),
    .gather_data_i                                     (gather_data_nw_2_pe[6][15]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[6][15]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[6][15]),
    .gather_data_o                                     (gather_data_pe_2_nw[6][15]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[6][15]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[6][15])
);


virtual_pe #(
    .cast_out                                          (cast_out_6_16),
    .merge_in                                          (merge_in_6_16),
    .merge_out                                         (merge_out_6_16),
    .gather_in                                         (gather_in_6_16),
    .gather_out                                        (gather_out_6_16),
    .x                                                 (6),
    .y                                                 (16)
)vpe_6_16(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[6][16]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[6][16]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[6][16]),
    .cast_data_o                                       (cast_data_pe_2_nw[6][16]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[6][16]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[6][16]),
    .merge_data_i                                      (merge_data_nw_2_pe[6][16]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[6][16]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[6][16]),
    .merge_data_o                                      (merge_data_pe_2_nw[6][16]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[6][16]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[6][16]),
    .gather_data_i                                     (gather_data_nw_2_pe[6][16]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[6][16]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[6][16]),
    .gather_data_o                                     (gather_data_pe_2_nw[6][16]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[6][16]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[6][16])
);


virtual_pe #(
    .cast_out                                          (cast_out_6_17),
    .merge_in                                          (merge_in_6_17),
    .merge_out                                         (merge_out_6_17),
    .gather_in                                         (gather_in_6_17),
    .gather_out                                        (gather_out_6_17),
    .x                                                 (6),
    .y                                                 (17)
)vpe_6_17(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[6][17]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[6][17]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[6][17]),
    .cast_data_o                                       (cast_data_pe_2_nw[6][17]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[6][17]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[6][17]),
    .merge_data_i                                      (merge_data_nw_2_pe[6][17]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[6][17]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[6][17]),
    .merge_data_o                                      (merge_data_pe_2_nw[6][17]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[6][17]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[6][17]),
    .gather_data_i                                     (gather_data_nw_2_pe[6][17]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[6][17]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[6][17]),
    .gather_data_o                                     (gather_data_pe_2_nw[6][17]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[6][17]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[6][17])
);


virtual_pe #(
    .cast_out                                          (cast_out_6_18),
    .merge_in                                          (merge_in_6_18),
    .merge_out                                         (merge_out_6_18),
    .gather_in                                         (gather_in_6_18),
    .gather_out                                        (gather_out_6_18),
    .x                                                 (6),
    .y                                                 (18)
)vpe_6_18(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[6][18]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[6][18]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[6][18]),
    .cast_data_o                                       (cast_data_pe_2_nw[6][18]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[6][18]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[6][18]),
    .merge_data_i                                      (merge_data_nw_2_pe[6][18]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[6][18]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[6][18]),
    .merge_data_o                                      (merge_data_pe_2_nw[6][18]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[6][18]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[6][18]),
    .gather_data_i                                     (gather_data_nw_2_pe[6][18]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[6][18]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[6][18]),
    .gather_data_o                                     (gather_data_pe_2_nw[6][18]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[6][18]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[6][18])
);


virtual_pe #(
    .cast_out                                          (cast_out_6_19),
    .merge_in                                          (merge_in_6_19),
    .merge_out                                         (merge_out_6_19),
    .gather_in                                         (gather_in_6_19),
    .gather_out                                        (gather_out_6_19),
    .x                                                 (6),
    .y                                                 (19)
)vpe_6_19(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[6][19]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[6][19]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[6][19]),
    .cast_data_o                                       (cast_data_pe_2_nw[6][19]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[6][19]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[6][19]),
    .merge_data_i                                      (merge_data_nw_2_pe[6][19]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[6][19]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[6][19]),
    .merge_data_o                                      (merge_data_pe_2_nw[6][19]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[6][19]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[6][19]),
    .gather_data_i                                     (gather_data_nw_2_pe[6][19]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[6][19]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[6][19]),
    .gather_data_o                                     (gather_data_pe_2_nw[6][19]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[6][19]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[6][19])
);


virtual_pe #(
    .cast_out                                          (cast_out_6_20),
    .merge_in                                          (merge_in_6_20),
    .merge_out                                         (merge_out_6_20),
    .gather_in                                         (gather_in_6_20),
    .gather_out                                        (gather_out_6_20),
    .x                                                 (6),
    .y                                                 (20)
)vpe_6_20(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[6][20]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[6][20]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[6][20]),
    .cast_data_o                                       (cast_data_pe_2_nw[6][20]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[6][20]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[6][20]),
    .merge_data_i                                      (merge_data_nw_2_pe[6][20]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[6][20]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[6][20]),
    .merge_data_o                                      (merge_data_pe_2_nw[6][20]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[6][20]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[6][20]),
    .gather_data_i                                     (gather_data_nw_2_pe[6][20]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[6][20]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[6][20]),
    .gather_data_o                                     (gather_data_pe_2_nw[6][20]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[6][20]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[6][20])
);


virtual_pe #(
    .cast_out                                          (cast_out_6_21),
    .merge_in                                          (merge_in_6_21),
    .merge_out                                         (merge_out_6_21),
    .gather_in                                         (gather_in_6_21),
    .gather_out                                        (gather_out_6_21),
    .x                                                 (6),
    .y                                                 (21)
)vpe_6_21(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[6][21]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[6][21]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[6][21]),
    .cast_data_o                                       (cast_data_pe_2_nw[6][21]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[6][21]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[6][21]),
    .merge_data_i                                      (merge_data_nw_2_pe[6][21]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[6][21]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[6][21]),
    .merge_data_o                                      (merge_data_pe_2_nw[6][21]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[6][21]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[6][21]),
    .gather_data_i                                     (gather_data_nw_2_pe[6][21]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[6][21]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[6][21]),
    .gather_data_o                                     (gather_data_pe_2_nw[6][21]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[6][21]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[6][21])
);


virtual_pe #(
    .cast_out                                          (cast_out_6_22),
    .merge_in                                          (merge_in_6_22),
    .merge_out                                         (merge_out_6_22),
    .gather_in                                         (gather_in_6_22),
    .gather_out                                        (gather_out_6_22),
    .x                                                 (6),
    .y                                                 (22)
)vpe_6_22(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[6][22]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[6][22]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[6][22]),
    .cast_data_o                                       (cast_data_pe_2_nw[6][22]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[6][22]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[6][22]),
    .merge_data_i                                      (merge_data_nw_2_pe[6][22]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[6][22]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[6][22]),
    .merge_data_o                                      (merge_data_pe_2_nw[6][22]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[6][22]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[6][22]),
    .gather_data_i                                     (gather_data_nw_2_pe[6][22]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[6][22]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[6][22]),
    .gather_data_o                                     (gather_data_pe_2_nw[6][22]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[6][22]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[6][22])
);


virtual_pe #(
    .cast_out                                          (cast_out_6_23),
    .merge_in                                          (merge_in_6_23),
    .merge_out                                         (merge_out_6_23),
    .gather_in                                         (gather_in_6_23),
    .gather_out                                        (gather_out_6_23),
    .x                                                 (6),
    .y                                                 (23)
)vpe_6_23(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[6][23]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[6][23]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[6][23]),
    .cast_data_o                                       (cast_data_pe_2_nw[6][23]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[6][23]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[6][23]),
    .merge_data_i                                      (merge_data_nw_2_pe[6][23]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[6][23]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[6][23]),
    .merge_data_o                                      (merge_data_pe_2_nw[6][23]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[6][23]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[6][23]),
    .gather_data_i                                     (gather_data_nw_2_pe[6][23]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[6][23]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[6][23]),
    .gather_data_o                                     (gather_data_pe_2_nw[6][23]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[6][23]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[6][23])
);


virtual_pe #(
    .cast_out                                          (cast_out_6_24),
    .merge_in                                          (merge_in_6_24),
    .merge_out                                         (merge_out_6_24),
    .gather_in                                         (gather_in_6_24),
    .gather_out                                        (gather_out_6_24),
    .x                                                 (6),
    .y                                                 (24)
)vpe_6_24(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[6][24]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[6][24]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[6][24]),
    .cast_data_o                                       (cast_data_pe_2_nw[6][24]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[6][24]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[6][24]),
    .merge_data_i                                      (merge_data_nw_2_pe[6][24]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[6][24]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[6][24]),
    .merge_data_o                                      (merge_data_pe_2_nw[6][24]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[6][24]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[6][24]),
    .gather_data_i                                     (gather_data_nw_2_pe[6][24]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[6][24]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[6][24]),
    .gather_data_o                                     (gather_data_pe_2_nw[6][24]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[6][24]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[6][24])
);


virtual_pe #(
    .cast_out                                          (cast_out_7_0),
    .merge_in                                          (merge_in_7_0),
    .merge_out                                         (merge_out_7_0),
    .gather_in                                         (gather_in_7_0),
    .gather_out                                        (gather_out_7_0),
    .x                                                 (7),
    .y                                                 (0)
)vpe_7_0(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[7][0]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[7][0]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[7][0]),
    .cast_data_o                                       (cast_data_pe_2_nw[7][0]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[7][0]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[7][0]),
    .merge_data_i                                      (merge_data_nw_2_pe[7][0]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[7][0]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[7][0]),
    .merge_data_o                                      (merge_data_pe_2_nw[7][0]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[7][0]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[7][0]),
    .gather_data_i                                     (gather_data_nw_2_pe[7][0]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[7][0]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[7][0]),
    .gather_data_o                                     (gather_data_pe_2_nw[7][0]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[7][0]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[7][0])
);


virtual_pe #(
    .cast_out                                          (cast_out_7_1),
    .merge_in                                          (merge_in_7_1),
    .merge_out                                         (merge_out_7_1),
    .gather_in                                         (gather_in_7_1),
    .gather_out                                        (gather_out_7_1),
    .x                                                 (7),
    .y                                                 (1)
)vpe_7_1(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[7][1]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[7][1]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[7][1]),
    .cast_data_o                                       (cast_data_pe_2_nw[7][1]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[7][1]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[7][1]),
    .merge_data_i                                      (merge_data_nw_2_pe[7][1]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[7][1]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[7][1]),
    .merge_data_o                                      (merge_data_pe_2_nw[7][1]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[7][1]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[7][1]),
    .gather_data_i                                     (gather_data_nw_2_pe[7][1]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[7][1]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[7][1]),
    .gather_data_o                                     (gather_data_pe_2_nw[7][1]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[7][1]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[7][1])
);


virtual_pe #(
    .cast_out                                          (cast_out_7_2),
    .merge_in                                          (merge_in_7_2),
    .merge_out                                         (merge_out_7_2),
    .gather_in                                         (gather_in_7_2),
    .gather_out                                        (gather_out_7_2),
    .x                                                 (7),
    .y                                                 (2)
)vpe_7_2(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[7][2]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[7][2]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[7][2]),
    .cast_data_o                                       (cast_data_pe_2_nw[7][2]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[7][2]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[7][2]),
    .merge_data_i                                      (merge_data_nw_2_pe[7][2]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[7][2]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[7][2]),
    .merge_data_o                                      (merge_data_pe_2_nw[7][2]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[7][2]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[7][2]),
    .gather_data_i                                     (gather_data_nw_2_pe[7][2]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[7][2]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[7][2]),
    .gather_data_o                                     (gather_data_pe_2_nw[7][2]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[7][2]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[7][2])
);


virtual_pe #(
    .cast_out                                          (cast_out_7_3),
    .merge_in                                          (merge_in_7_3),
    .merge_out                                         (merge_out_7_3),
    .gather_in                                         (gather_in_7_3),
    .gather_out                                        (gather_out_7_3),
    .x                                                 (7),
    .y                                                 (3)
)vpe_7_3(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[7][3]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[7][3]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[7][3]),
    .cast_data_o                                       (cast_data_pe_2_nw[7][3]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[7][3]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[7][3]),
    .merge_data_i                                      (merge_data_nw_2_pe[7][3]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[7][3]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[7][3]),
    .merge_data_o                                      (merge_data_pe_2_nw[7][3]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[7][3]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[7][3]),
    .gather_data_i                                     (gather_data_nw_2_pe[7][3]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[7][3]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[7][3]),
    .gather_data_o                                     (gather_data_pe_2_nw[7][3]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[7][3]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[7][3])
);


virtual_pe #(
    .cast_out                                          (cast_out_7_4),
    .merge_in                                          (merge_in_7_4),
    .merge_out                                         (merge_out_7_4),
    .gather_in                                         (gather_in_7_4),
    .gather_out                                        (gather_out_7_4),
    .x                                                 (7),
    .y                                                 (4)
)vpe_7_4(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[7][4]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[7][4]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[7][4]),
    .cast_data_o                                       (cast_data_pe_2_nw[7][4]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[7][4]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[7][4]),
    .merge_data_i                                      (merge_data_nw_2_pe[7][4]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[7][4]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[7][4]),
    .merge_data_o                                      (merge_data_pe_2_nw[7][4]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[7][4]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[7][4]),
    .gather_data_i                                     (gather_data_nw_2_pe[7][4]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[7][4]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[7][4]),
    .gather_data_o                                     (gather_data_pe_2_nw[7][4]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[7][4]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[7][4])
);


virtual_pe #(
    .cast_out                                          (cast_out_7_5),
    .merge_in                                          (merge_in_7_5),
    .merge_out                                         (merge_out_7_5),
    .gather_in                                         (gather_in_7_5),
    .gather_out                                        (gather_out_7_5),
    .x                                                 (7),
    .y                                                 (5)
)vpe_7_5(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[7][5]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[7][5]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[7][5]),
    .cast_data_o                                       (cast_data_pe_2_nw[7][5]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[7][5]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[7][5]),
    .merge_data_i                                      (merge_data_nw_2_pe[7][5]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[7][5]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[7][5]),
    .merge_data_o                                      (merge_data_pe_2_nw[7][5]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[7][5]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[7][5]),
    .gather_data_i                                     (gather_data_nw_2_pe[7][5]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[7][5]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[7][5]),
    .gather_data_o                                     (gather_data_pe_2_nw[7][5]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[7][5]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[7][5])
);


virtual_pe #(
    .cast_out                                          (cast_out_7_6),
    .merge_in                                          (merge_in_7_6),
    .merge_out                                         (merge_out_7_6),
    .gather_in                                         (gather_in_7_6),
    .gather_out                                        (gather_out_7_6),
    .x                                                 (7),
    .y                                                 (6)
)vpe_7_6(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[7][6]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[7][6]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[7][6]),
    .cast_data_o                                       (cast_data_pe_2_nw[7][6]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[7][6]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[7][6]),
    .merge_data_i                                      (merge_data_nw_2_pe[7][6]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[7][6]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[7][6]),
    .merge_data_o                                      (merge_data_pe_2_nw[7][6]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[7][6]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[7][6]),
    .gather_data_i                                     (gather_data_nw_2_pe[7][6]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[7][6]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[7][6]),
    .gather_data_o                                     (gather_data_pe_2_nw[7][6]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[7][6]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[7][6])
);


virtual_pe #(
    .cast_out                                          (cast_out_7_7),
    .merge_in                                          (merge_in_7_7),
    .merge_out                                         (merge_out_7_7),
    .gather_in                                         (gather_in_7_7),
    .gather_out                                        (gather_out_7_7),
    .x                                                 (7),
    .y                                                 (7)
)vpe_7_7(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[7][7]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[7][7]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[7][7]),
    .cast_data_o                                       (cast_data_pe_2_nw[7][7]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[7][7]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[7][7]),
    .merge_data_i                                      (merge_data_nw_2_pe[7][7]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[7][7]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[7][7]),
    .merge_data_o                                      (merge_data_pe_2_nw[7][7]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[7][7]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[7][7]),
    .gather_data_i                                     (gather_data_nw_2_pe[7][7]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[7][7]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[7][7]),
    .gather_data_o                                     (gather_data_pe_2_nw[7][7]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[7][7]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[7][7])
);


virtual_pe #(
    .cast_out                                          (cast_out_7_8),
    .merge_in                                          (merge_in_7_8),
    .merge_out                                         (merge_out_7_8),
    .gather_in                                         (gather_in_7_8),
    .gather_out                                        (gather_out_7_8),
    .x                                                 (7),
    .y                                                 (8)
)vpe_7_8(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[7][8]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[7][8]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[7][8]),
    .cast_data_o                                       (cast_data_pe_2_nw[7][8]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[7][8]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[7][8]),
    .merge_data_i                                      (merge_data_nw_2_pe[7][8]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[7][8]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[7][8]),
    .merge_data_o                                      (merge_data_pe_2_nw[7][8]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[7][8]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[7][8]),
    .gather_data_i                                     (gather_data_nw_2_pe[7][8]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[7][8]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[7][8]),
    .gather_data_o                                     (gather_data_pe_2_nw[7][8]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[7][8]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[7][8])
);


virtual_pe #(
    .cast_out                                          (cast_out_7_9),
    .merge_in                                          (merge_in_7_9),
    .merge_out                                         (merge_out_7_9),
    .gather_in                                         (gather_in_7_9),
    .gather_out                                        (gather_out_7_9),
    .x                                                 (7),
    .y                                                 (9)
)vpe_7_9(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[7][9]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[7][9]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[7][9]),
    .cast_data_o                                       (cast_data_pe_2_nw[7][9]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[7][9]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[7][9]),
    .merge_data_i                                      (merge_data_nw_2_pe[7][9]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[7][9]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[7][9]),
    .merge_data_o                                      (merge_data_pe_2_nw[7][9]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[7][9]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[7][9]),
    .gather_data_i                                     (gather_data_nw_2_pe[7][9]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[7][9]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[7][9]),
    .gather_data_o                                     (gather_data_pe_2_nw[7][9]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[7][9]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[7][9])
);


virtual_pe #(
    .cast_out                                          (cast_out_7_10),
    .merge_in                                          (merge_in_7_10),
    .merge_out                                         (merge_out_7_10),
    .gather_in                                         (gather_in_7_10),
    .gather_out                                        (gather_out_7_10),
    .x                                                 (7),
    .y                                                 (10)
)vpe_7_10(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[7][10]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[7][10]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[7][10]),
    .cast_data_o                                       (cast_data_pe_2_nw[7][10]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[7][10]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[7][10]),
    .merge_data_i                                      (merge_data_nw_2_pe[7][10]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[7][10]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[7][10]),
    .merge_data_o                                      (merge_data_pe_2_nw[7][10]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[7][10]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[7][10]),
    .gather_data_i                                     (gather_data_nw_2_pe[7][10]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[7][10]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[7][10]),
    .gather_data_o                                     (gather_data_pe_2_nw[7][10]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[7][10]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[7][10])
);


virtual_pe #(
    .cast_out                                          (cast_out_7_11),
    .merge_in                                          (merge_in_7_11),
    .merge_out                                         (merge_out_7_11),
    .gather_in                                         (gather_in_7_11),
    .gather_out                                        (gather_out_7_11),
    .x                                                 (7),
    .y                                                 (11)
)vpe_7_11(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[7][11]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[7][11]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[7][11]),
    .cast_data_o                                       (cast_data_pe_2_nw[7][11]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[7][11]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[7][11]),
    .merge_data_i                                      (merge_data_nw_2_pe[7][11]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[7][11]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[7][11]),
    .merge_data_o                                      (merge_data_pe_2_nw[7][11]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[7][11]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[7][11]),
    .gather_data_i                                     (gather_data_nw_2_pe[7][11]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[7][11]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[7][11]),
    .gather_data_o                                     (gather_data_pe_2_nw[7][11]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[7][11]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[7][11])
);


virtual_pe #(
    .cast_out                                          (cast_out_7_12),
    .merge_in                                          (merge_in_7_12),
    .merge_out                                         (merge_out_7_12),
    .gather_in                                         (gather_in_7_12),
    .gather_out                                        (gather_out_7_12),
    .x                                                 (7),
    .y                                                 (12)
)vpe_7_12(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[7][12]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[7][12]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[7][12]),
    .cast_data_o                                       (cast_data_pe_2_nw[7][12]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[7][12]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[7][12]),
    .merge_data_i                                      (merge_data_nw_2_pe[7][12]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[7][12]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[7][12]),
    .merge_data_o                                      (merge_data_pe_2_nw[7][12]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[7][12]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[7][12]),
    .gather_data_i                                     (gather_data_nw_2_pe[7][12]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[7][12]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[7][12]),
    .gather_data_o                                     (gather_data_pe_2_nw[7][12]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[7][12]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[7][12])
);


virtual_pe #(
    .cast_out                                          (cast_out_7_13),
    .merge_in                                          (merge_in_7_13),
    .merge_out                                         (merge_out_7_13),
    .gather_in                                         (gather_in_7_13),
    .gather_out                                        (gather_out_7_13),
    .x                                                 (7),
    .y                                                 (13)
)vpe_7_13(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[7][13]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[7][13]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[7][13]),
    .cast_data_o                                       (cast_data_pe_2_nw[7][13]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[7][13]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[7][13]),
    .merge_data_i                                      (merge_data_nw_2_pe[7][13]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[7][13]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[7][13]),
    .merge_data_o                                      (merge_data_pe_2_nw[7][13]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[7][13]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[7][13]),
    .gather_data_i                                     (gather_data_nw_2_pe[7][13]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[7][13]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[7][13]),
    .gather_data_o                                     (gather_data_pe_2_nw[7][13]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[7][13]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[7][13])
);


virtual_pe #(
    .cast_out                                          (cast_out_7_14),
    .merge_in                                          (merge_in_7_14),
    .merge_out                                         (merge_out_7_14),
    .gather_in                                         (gather_in_7_14),
    .gather_out                                        (gather_out_7_14),
    .x                                                 (7),
    .y                                                 (14)
)vpe_7_14(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[7][14]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[7][14]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[7][14]),
    .cast_data_o                                       (cast_data_pe_2_nw[7][14]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[7][14]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[7][14]),
    .merge_data_i                                      (merge_data_nw_2_pe[7][14]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[7][14]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[7][14]),
    .merge_data_o                                      (merge_data_pe_2_nw[7][14]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[7][14]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[7][14]),
    .gather_data_i                                     (gather_data_nw_2_pe[7][14]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[7][14]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[7][14]),
    .gather_data_o                                     (gather_data_pe_2_nw[7][14]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[7][14]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[7][14])
);


virtual_pe #(
    .cast_out                                          (cast_out_7_15),
    .merge_in                                          (merge_in_7_15),
    .merge_out                                         (merge_out_7_15),
    .gather_in                                         (gather_in_7_15),
    .gather_out                                        (gather_out_7_15),
    .x                                                 (7),
    .y                                                 (15)
)vpe_7_15(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[7][15]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[7][15]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[7][15]),
    .cast_data_o                                       (cast_data_pe_2_nw[7][15]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[7][15]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[7][15]),
    .merge_data_i                                      (merge_data_nw_2_pe[7][15]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[7][15]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[7][15]),
    .merge_data_o                                      (merge_data_pe_2_nw[7][15]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[7][15]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[7][15]),
    .gather_data_i                                     (gather_data_nw_2_pe[7][15]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[7][15]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[7][15]),
    .gather_data_o                                     (gather_data_pe_2_nw[7][15]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[7][15]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[7][15])
);


virtual_pe #(
    .cast_out                                          (cast_out_7_16),
    .merge_in                                          (merge_in_7_16),
    .merge_out                                         (merge_out_7_16),
    .gather_in                                         (gather_in_7_16),
    .gather_out                                        (gather_out_7_16),
    .x                                                 (7),
    .y                                                 (16)
)vpe_7_16(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[7][16]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[7][16]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[7][16]),
    .cast_data_o                                       (cast_data_pe_2_nw[7][16]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[7][16]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[7][16]),
    .merge_data_i                                      (merge_data_nw_2_pe[7][16]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[7][16]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[7][16]),
    .merge_data_o                                      (merge_data_pe_2_nw[7][16]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[7][16]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[7][16]),
    .gather_data_i                                     (gather_data_nw_2_pe[7][16]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[7][16]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[7][16]),
    .gather_data_o                                     (gather_data_pe_2_nw[7][16]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[7][16]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[7][16])
);


virtual_pe #(
    .cast_out                                          (cast_out_7_17),
    .merge_in                                          (merge_in_7_17),
    .merge_out                                         (merge_out_7_17),
    .gather_in                                         (gather_in_7_17),
    .gather_out                                        (gather_out_7_17),
    .x                                                 (7),
    .y                                                 (17)
)vpe_7_17(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[7][17]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[7][17]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[7][17]),
    .cast_data_o                                       (cast_data_pe_2_nw[7][17]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[7][17]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[7][17]),
    .merge_data_i                                      (merge_data_nw_2_pe[7][17]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[7][17]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[7][17]),
    .merge_data_o                                      (merge_data_pe_2_nw[7][17]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[7][17]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[7][17]),
    .gather_data_i                                     (gather_data_nw_2_pe[7][17]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[7][17]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[7][17]),
    .gather_data_o                                     (gather_data_pe_2_nw[7][17]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[7][17]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[7][17])
);


virtual_pe #(
    .cast_out                                          (cast_out_7_18),
    .merge_in                                          (merge_in_7_18),
    .merge_out                                         (merge_out_7_18),
    .gather_in                                         (gather_in_7_18),
    .gather_out                                        (gather_out_7_18),
    .x                                                 (7),
    .y                                                 (18)
)vpe_7_18(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[7][18]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[7][18]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[7][18]),
    .cast_data_o                                       (cast_data_pe_2_nw[7][18]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[7][18]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[7][18]),
    .merge_data_i                                      (merge_data_nw_2_pe[7][18]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[7][18]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[7][18]),
    .merge_data_o                                      (merge_data_pe_2_nw[7][18]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[7][18]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[7][18]),
    .gather_data_i                                     (gather_data_nw_2_pe[7][18]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[7][18]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[7][18]),
    .gather_data_o                                     (gather_data_pe_2_nw[7][18]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[7][18]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[7][18])
);


virtual_pe #(
    .cast_out                                          (cast_out_7_19),
    .merge_in                                          (merge_in_7_19),
    .merge_out                                         (merge_out_7_19),
    .gather_in                                         (gather_in_7_19),
    .gather_out                                        (gather_out_7_19),
    .x                                                 (7),
    .y                                                 (19)
)vpe_7_19(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[7][19]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[7][19]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[7][19]),
    .cast_data_o                                       (cast_data_pe_2_nw[7][19]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[7][19]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[7][19]),
    .merge_data_i                                      (merge_data_nw_2_pe[7][19]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[7][19]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[7][19]),
    .merge_data_o                                      (merge_data_pe_2_nw[7][19]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[7][19]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[7][19]),
    .gather_data_i                                     (gather_data_nw_2_pe[7][19]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[7][19]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[7][19]),
    .gather_data_o                                     (gather_data_pe_2_nw[7][19]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[7][19]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[7][19])
);


virtual_pe #(
    .cast_out                                          (cast_out_7_20),
    .merge_in                                          (merge_in_7_20),
    .merge_out                                         (merge_out_7_20),
    .gather_in                                         (gather_in_7_20),
    .gather_out                                        (gather_out_7_20),
    .x                                                 (7),
    .y                                                 (20)
)vpe_7_20(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[7][20]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[7][20]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[7][20]),
    .cast_data_o                                       (cast_data_pe_2_nw[7][20]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[7][20]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[7][20]),
    .merge_data_i                                      (merge_data_nw_2_pe[7][20]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[7][20]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[7][20]),
    .merge_data_o                                      (merge_data_pe_2_nw[7][20]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[7][20]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[7][20]),
    .gather_data_i                                     (gather_data_nw_2_pe[7][20]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[7][20]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[7][20]),
    .gather_data_o                                     (gather_data_pe_2_nw[7][20]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[7][20]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[7][20])
);


virtual_pe #(
    .cast_out                                          (cast_out_7_21),
    .merge_in                                          (merge_in_7_21),
    .merge_out                                         (merge_out_7_21),
    .gather_in                                         (gather_in_7_21),
    .gather_out                                        (gather_out_7_21),
    .x                                                 (7),
    .y                                                 (21)
)vpe_7_21(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[7][21]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[7][21]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[7][21]),
    .cast_data_o                                       (cast_data_pe_2_nw[7][21]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[7][21]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[7][21]),
    .merge_data_i                                      (merge_data_nw_2_pe[7][21]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[7][21]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[7][21]),
    .merge_data_o                                      (merge_data_pe_2_nw[7][21]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[7][21]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[7][21]),
    .gather_data_i                                     (gather_data_nw_2_pe[7][21]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[7][21]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[7][21]),
    .gather_data_o                                     (gather_data_pe_2_nw[7][21]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[7][21]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[7][21])
);


virtual_pe #(
    .cast_out                                          (cast_out_7_22),
    .merge_in                                          (merge_in_7_22),
    .merge_out                                         (merge_out_7_22),
    .gather_in                                         (gather_in_7_22),
    .gather_out                                        (gather_out_7_22),
    .x                                                 (7),
    .y                                                 (22)
)vpe_7_22(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[7][22]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[7][22]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[7][22]),
    .cast_data_o                                       (cast_data_pe_2_nw[7][22]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[7][22]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[7][22]),
    .merge_data_i                                      (merge_data_nw_2_pe[7][22]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[7][22]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[7][22]),
    .merge_data_o                                      (merge_data_pe_2_nw[7][22]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[7][22]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[7][22]),
    .gather_data_i                                     (gather_data_nw_2_pe[7][22]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[7][22]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[7][22]),
    .gather_data_o                                     (gather_data_pe_2_nw[7][22]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[7][22]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[7][22])
);


virtual_pe #(
    .cast_out                                          (cast_out_7_23),
    .merge_in                                          (merge_in_7_23),
    .merge_out                                         (merge_out_7_23),
    .gather_in                                         (gather_in_7_23),
    .gather_out                                        (gather_out_7_23),
    .x                                                 (7),
    .y                                                 (23)
)vpe_7_23(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[7][23]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[7][23]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[7][23]),
    .cast_data_o                                       (cast_data_pe_2_nw[7][23]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[7][23]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[7][23]),
    .merge_data_i                                      (merge_data_nw_2_pe[7][23]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[7][23]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[7][23]),
    .merge_data_o                                      (merge_data_pe_2_nw[7][23]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[7][23]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[7][23]),
    .gather_data_i                                     (gather_data_nw_2_pe[7][23]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[7][23]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[7][23]),
    .gather_data_o                                     (gather_data_pe_2_nw[7][23]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[7][23]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[7][23])
);


virtual_pe #(
    .cast_out                                          (cast_out_7_24),
    .merge_in                                          (merge_in_7_24),
    .merge_out                                         (merge_out_7_24),
    .gather_in                                         (gather_in_7_24),
    .gather_out                                        (gather_out_7_24),
    .x                                                 (7),
    .y                                                 (24)
)vpe_7_24(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[7][24]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[7][24]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[7][24]),
    .cast_data_o                                       (cast_data_pe_2_nw[7][24]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[7][24]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[7][24]),
    .merge_data_i                                      (merge_data_nw_2_pe[7][24]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[7][24]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[7][24]),
    .merge_data_o                                      (merge_data_pe_2_nw[7][24]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[7][24]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[7][24]),
    .gather_data_i                                     (gather_data_nw_2_pe[7][24]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[7][24]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[7][24]),
    .gather_data_o                                     (gather_data_pe_2_nw[7][24]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[7][24]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[7][24])
);


virtual_pe #(
    .cast_out                                          (cast_out_8_0),
    .merge_in                                          (merge_in_8_0),
    .merge_out                                         (merge_out_8_0),
    .gather_in                                         (gather_in_8_0),
    .gather_out                                        (gather_out_8_0),
    .x                                                 (8),
    .y                                                 (0)
)vpe_8_0(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[8][0]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[8][0]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[8][0]),
    .cast_data_o                                       (cast_data_pe_2_nw[8][0]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[8][0]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[8][0]),
    .merge_data_i                                      (merge_data_nw_2_pe[8][0]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[8][0]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[8][0]),
    .merge_data_o                                      (merge_data_pe_2_nw[8][0]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[8][0]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[8][0]),
    .gather_data_i                                     (gather_data_nw_2_pe[8][0]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[8][0]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[8][0]),
    .gather_data_o                                     (gather_data_pe_2_nw[8][0]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[8][0]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[8][0])
);


virtual_pe #(
    .cast_out                                          (cast_out_8_1),
    .merge_in                                          (merge_in_8_1),
    .merge_out                                         (merge_out_8_1),
    .gather_in                                         (gather_in_8_1),
    .gather_out                                        (gather_out_8_1),
    .x                                                 (8),
    .y                                                 (1)
)vpe_8_1(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[8][1]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[8][1]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[8][1]),
    .cast_data_o                                       (cast_data_pe_2_nw[8][1]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[8][1]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[8][1]),
    .merge_data_i                                      (merge_data_nw_2_pe[8][1]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[8][1]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[8][1]),
    .merge_data_o                                      (merge_data_pe_2_nw[8][1]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[8][1]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[8][1]),
    .gather_data_i                                     (gather_data_nw_2_pe[8][1]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[8][1]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[8][1]),
    .gather_data_o                                     (gather_data_pe_2_nw[8][1]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[8][1]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[8][1])
);


virtual_pe #(
    .cast_out                                          (cast_out_8_2),
    .merge_in                                          (merge_in_8_2),
    .merge_out                                         (merge_out_8_2),
    .gather_in                                         (gather_in_8_2),
    .gather_out                                        (gather_out_8_2),
    .x                                                 (8),
    .y                                                 (2)
)vpe_8_2(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[8][2]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[8][2]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[8][2]),
    .cast_data_o                                       (cast_data_pe_2_nw[8][2]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[8][2]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[8][2]),
    .merge_data_i                                      (merge_data_nw_2_pe[8][2]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[8][2]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[8][2]),
    .merge_data_o                                      (merge_data_pe_2_nw[8][2]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[8][2]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[8][2]),
    .gather_data_i                                     (gather_data_nw_2_pe[8][2]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[8][2]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[8][2]),
    .gather_data_o                                     (gather_data_pe_2_nw[8][2]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[8][2]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[8][2])
);


virtual_pe #(
    .cast_out                                          (cast_out_8_3),
    .merge_in                                          (merge_in_8_3),
    .merge_out                                         (merge_out_8_3),
    .gather_in                                         (gather_in_8_3),
    .gather_out                                        (gather_out_8_3),
    .x                                                 (8),
    .y                                                 (3)
)vpe_8_3(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[8][3]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[8][3]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[8][3]),
    .cast_data_o                                       (cast_data_pe_2_nw[8][3]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[8][3]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[8][3]),
    .merge_data_i                                      (merge_data_nw_2_pe[8][3]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[8][3]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[8][3]),
    .merge_data_o                                      (merge_data_pe_2_nw[8][3]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[8][3]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[8][3]),
    .gather_data_i                                     (gather_data_nw_2_pe[8][3]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[8][3]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[8][3]),
    .gather_data_o                                     (gather_data_pe_2_nw[8][3]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[8][3]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[8][3])
);


virtual_pe #(
    .cast_out                                          (cast_out_8_4),
    .merge_in                                          (merge_in_8_4),
    .merge_out                                         (merge_out_8_4),
    .gather_in                                         (gather_in_8_4),
    .gather_out                                        (gather_out_8_4),
    .x                                                 (8),
    .y                                                 (4)
)vpe_8_4(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[8][4]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[8][4]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[8][4]),
    .cast_data_o                                       (cast_data_pe_2_nw[8][4]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[8][4]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[8][4]),
    .merge_data_i                                      (merge_data_nw_2_pe[8][4]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[8][4]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[8][4]),
    .merge_data_o                                      (merge_data_pe_2_nw[8][4]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[8][4]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[8][4]),
    .gather_data_i                                     (gather_data_nw_2_pe[8][4]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[8][4]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[8][4]),
    .gather_data_o                                     (gather_data_pe_2_nw[8][4]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[8][4]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[8][4])
);


virtual_pe #(
    .cast_out                                          (cast_out_8_5),
    .merge_in                                          (merge_in_8_5),
    .merge_out                                         (merge_out_8_5),
    .gather_in                                         (gather_in_8_5),
    .gather_out                                        (gather_out_8_5),
    .x                                                 (8),
    .y                                                 (5)
)vpe_8_5(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[8][5]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[8][5]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[8][5]),
    .cast_data_o                                       (cast_data_pe_2_nw[8][5]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[8][5]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[8][5]),
    .merge_data_i                                      (merge_data_nw_2_pe[8][5]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[8][5]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[8][5]),
    .merge_data_o                                      (merge_data_pe_2_nw[8][5]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[8][5]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[8][5]),
    .gather_data_i                                     (gather_data_nw_2_pe[8][5]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[8][5]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[8][5]),
    .gather_data_o                                     (gather_data_pe_2_nw[8][5]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[8][5]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[8][5])
);


virtual_pe #(
    .cast_out                                          (cast_out_8_6),
    .merge_in                                          (merge_in_8_6),
    .merge_out                                         (merge_out_8_6),
    .gather_in                                         (gather_in_8_6),
    .gather_out                                        (gather_out_8_6),
    .x                                                 (8),
    .y                                                 (6)
)vpe_8_6(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[8][6]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[8][6]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[8][6]),
    .cast_data_o                                       (cast_data_pe_2_nw[8][6]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[8][6]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[8][6]),
    .merge_data_i                                      (merge_data_nw_2_pe[8][6]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[8][6]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[8][6]),
    .merge_data_o                                      (merge_data_pe_2_nw[8][6]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[8][6]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[8][6]),
    .gather_data_i                                     (gather_data_nw_2_pe[8][6]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[8][6]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[8][6]),
    .gather_data_o                                     (gather_data_pe_2_nw[8][6]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[8][6]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[8][6])
);


virtual_pe #(
    .cast_out                                          (cast_out_8_7),
    .merge_in                                          (merge_in_8_7),
    .merge_out                                         (merge_out_8_7),
    .gather_in                                         (gather_in_8_7),
    .gather_out                                        (gather_out_8_7),
    .x                                                 (8),
    .y                                                 (7)
)vpe_8_7(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[8][7]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[8][7]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[8][7]),
    .cast_data_o                                       (cast_data_pe_2_nw[8][7]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[8][7]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[8][7]),
    .merge_data_i                                      (merge_data_nw_2_pe[8][7]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[8][7]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[8][7]),
    .merge_data_o                                      (merge_data_pe_2_nw[8][7]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[8][7]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[8][7]),
    .gather_data_i                                     (gather_data_nw_2_pe[8][7]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[8][7]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[8][7]),
    .gather_data_o                                     (gather_data_pe_2_nw[8][7]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[8][7]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[8][7])
);


virtual_pe #(
    .cast_out                                          (cast_out_8_8),
    .merge_in                                          (merge_in_8_8),
    .merge_out                                         (merge_out_8_8),
    .gather_in                                         (gather_in_8_8),
    .gather_out                                        (gather_out_8_8),
    .x                                                 (8),
    .y                                                 (8)
)vpe_8_8(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[8][8]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[8][8]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[8][8]),
    .cast_data_o                                       (cast_data_pe_2_nw[8][8]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[8][8]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[8][8]),
    .merge_data_i                                      (merge_data_nw_2_pe[8][8]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[8][8]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[8][8]),
    .merge_data_o                                      (merge_data_pe_2_nw[8][8]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[8][8]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[8][8]),
    .gather_data_i                                     (gather_data_nw_2_pe[8][8]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[8][8]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[8][8]),
    .gather_data_o                                     (gather_data_pe_2_nw[8][8]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[8][8]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[8][8])
);


virtual_pe #(
    .cast_out                                          (cast_out_8_9),
    .merge_in                                          (merge_in_8_9),
    .merge_out                                         (merge_out_8_9),
    .gather_in                                         (gather_in_8_9),
    .gather_out                                        (gather_out_8_9),
    .x                                                 (8),
    .y                                                 (9)
)vpe_8_9(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[8][9]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[8][9]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[8][9]),
    .cast_data_o                                       (cast_data_pe_2_nw[8][9]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[8][9]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[8][9]),
    .merge_data_i                                      (merge_data_nw_2_pe[8][9]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[8][9]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[8][9]),
    .merge_data_o                                      (merge_data_pe_2_nw[8][9]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[8][9]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[8][9]),
    .gather_data_i                                     (gather_data_nw_2_pe[8][9]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[8][9]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[8][9]),
    .gather_data_o                                     (gather_data_pe_2_nw[8][9]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[8][9]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[8][9])
);


virtual_pe #(
    .cast_out                                          (cast_out_8_10),
    .merge_in                                          (merge_in_8_10),
    .merge_out                                         (merge_out_8_10),
    .gather_in                                         (gather_in_8_10),
    .gather_out                                        (gather_out_8_10),
    .x                                                 (8),
    .y                                                 (10)
)vpe_8_10(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[8][10]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[8][10]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[8][10]),
    .cast_data_o                                       (cast_data_pe_2_nw[8][10]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[8][10]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[8][10]),
    .merge_data_i                                      (merge_data_nw_2_pe[8][10]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[8][10]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[8][10]),
    .merge_data_o                                      (merge_data_pe_2_nw[8][10]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[8][10]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[8][10]),
    .gather_data_i                                     (gather_data_nw_2_pe[8][10]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[8][10]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[8][10]),
    .gather_data_o                                     (gather_data_pe_2_nw[8][10]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[8][10]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[8][10])
);


virtual_pe #(
    .cast_out                                          (cast_out_8_11),
    .merge_in                                          (merge_in_8_11),
    .merge_out                                         (merge_out_8_11),
    .gather_in                                         (gather_in_8_11),
    .gather_out                                        (gather_out_8_11),
    .x                                                 (8),
    .y                                                 (11)
)vpe_8_11(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[8][11]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[8][11]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[8][11]),
    .cast_data_o                                       (cast_data_pe_2_nw[8][11]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[8][11]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[8][11]),
    .merge_data_i                                      (merge_data_nw_2_pe[8][11]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[8][11]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[8][11]),
    .merge_data_o                                      (merge_data_pe_2_nw[8][11]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[8][11]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[8][11]),
    .gather_data_i                                     (gather_data_nw_2_pe[8][11]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[8][11]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[8][11]),
    .gather_data_o                                     (gather_data_pe_2_nw[8][11]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[8][11]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[8][11])
);


virtual_pe #(
    .cast_out                                          (cast_out_8_12),
    .merge_in                                          (merge_in_8_12),
    .merge_out                                         (merge_out_8_12),
    .gather_in                                         (gather_in_8_12),
    .gather_out                                        (gather_out_8_12),
    .x                                                 (8),
    .y                                                 (12)
)vpe_8_12(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[8][12]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[8][12]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[8][12]),
    .cast_data_o                                       (cast_data_pe_2_nw[8][12]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[8][12]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[8][12]),
    .merge_data_i                                      (merge_data_nw_2_pe[8][12]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[8][12]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[8][12]),
    .merge_data_o                                      (merge_data_pe_2_nw[8][12]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[8][12]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[8][12]),
    .gather_data_i                                     (gather_data_nw_2_pe[8][12]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[8][12]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[8][12]),
    .gather_data_o                                     (gather_data_pe_2_nw[8][12]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[8][12]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[8][12])
);


virtual_pe #(
    .cast_out                                          (cast_out_8_13),
    .merge_in                                          (merge_in_8_13),
    .merge_out                                         (merge_out_8_13),
    .gather_in                                         (gather_in_8_13),
    .gather_out                                        (gather_out_8_13),
    .x                                                 (8),
    .y                                                 (13)
)vpe_8_13(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[8][13]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[8][13]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[8][13]),
    .cast_data_o                                       (cast_data_pe_2_nw[8][13]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[8][13]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[8][13]),
    .merge_data_i                                      (merge_data_nw_2_pe[8][13]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[8][13]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[8][13]),
    .merge_data_o                                      (merge_data_pe_2_nw[8][13]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[8][13]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[8][13]),
    .gather_data_i                                     (gather_data_nw_2_pe[8][13]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[8][13]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[8][13]),
    .gather_data_o                                     (gather_data_pe_2_nw[8][13]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[8][13]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[8][13])
);


virtual_pe #(
    .cast_out                                          (cast_out_8_14),
    .merge_in                                          (merge_in_8_14),
    .merge_out                                         (merge_out_8_14),
    .gather_in                                         (gather_in_8_14),
    .gather_out                                        (gather_out_8_14),
    .x                                                 (8),
    .y                                                 (14)
)vpe_8_14(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[8][14]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[8][14]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[8][14]),
    .cast_data_o                                       (cast_data_pe_2_nw[8][14]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[8][14]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[8][14]),
    .merge_data_i                                      (merge_data_nw_2_pe[8][14]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[8][14]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[8][14]),
    .merge_data_o                                      (merge_data_pe_2_nw[8][14]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[8][14]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[8][14]),
    .gather_data_i                                     (gather_data_nw_2_pe[8][14]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[8][14]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[8][14]),
    .gather_data_o                                     (gather_data_pe_2_nw[8][14]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[8][14]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[8][14])
);


virtual_pe #(
    .cast_out                                          (cast_out_8_15),
    .merge_in                                          (merge_in_8_15),
    .merge_out                                         (merge_out_8_15),
    .gather_in                                         (gather_in_8_15),
    .gather_out                                        (gather_out_8_15),
    .x                                                 (8),
    .y                                                 (15)
)vpe_8_15(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[8][15]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[8][15]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[8][15]),
    .cast_data_o                                       (cast_data_pe_2_nw[8][15]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[8][15]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[8][15]),
    .merge_data_i                                      (merge_data_nw_2_pe[8][15]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[8][15]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[8][15]),
    .merge_data_o                                      (merge_data_pe_2_nw[8][15]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[8][15]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[8][15]),
    .gather_data_i                                     (gather_data_nw_2_pe[8][15]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[8][15]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[8][15]),
    .gather_data_o                                     (gather_data_pe_2_nw[8][15]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[8][15]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[8][15])
);


virtual_pe #(
    .cast_out                                          (cast_out_8_16),
    .merge_in                                          (merge_in_8_16),
    .merge_out                                         (merge_out_8_16),
    .gather_in                                         (gather_in_8_16),
    .gather_out                                        (gather_out_8_16),
    .x                                                 (8),
    .y                                                 (16)
)vpe_8_16(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[8][16]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[8][16]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[8][16]),
    .cast_data_o                                       (cast_data_pe_2_nw[8][16]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[8][16]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[8][16]),
    .merge_data_i                                      (merge_data_nw_2_pe[8][16]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[8][16]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[8][16]),
    .merge_data_o                                      (merge_data_pe_2_nw[8][16]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[8][16]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[8][16]),
    .gather_data_i                                     (gather_data_nw_2_pe[8][16]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[8][16]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[8][16]),
    .gather_data_o                                     (gather_data_pe_2_nw[8][16]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[8][16]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[8][16])
);


virtual_pe #(
    .cast_out                                          (cast_out_8_17),
    .merge_in                                          (merge_in_8_17),
    .merge_out                                         (merge_out_8_17),
    .gather_in                                         (gather_in_8_17),
    .gather_out                                        (gather_out_8_17),
    .x                                                 (8),
    .y                                                 (17)
)vpe_8_17(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[8][17]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[8][17]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[8][17]),
    .cast_data_o                                       (cast_data_pe_2_nw[8][17]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[8][17]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[8][17]),
    .merge_data_i                                      (merge_data_nw_2_pe[8][17]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[8][17]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[8][17]),
    .merge_data_o                                      (merge_data_pe_2_nw[8][17]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[8][17]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[8][17]),
    .gather_data_i                                     (gather_data_nw_2_pe[8][17]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[8][17]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[8][17]),
    .gather_data_o                                     (gather_data_pe_2_nw[8][17]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[8][17]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[8][17])
);


virtual_pe #(
    .cast_out                                          (cast_out_8_18),
    .merge_in                                          (merge_in_8_18),
    .merge_out                                         (merge_out_8_18),
    .gather_in                                         (gather_in_8_18),
    .gather_out                                        (gather_out_8_18),
    .x                                                 (8),
    .y                                                 (18)
)vpe_8_18(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[8][18]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[8][18]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[8][18]),
    .cast_data_o                                       (cast_data_pe_2_nw[8][18]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[8][18]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[8][18]),
    .merge_data_i                                      (merge_data_nw_2_pe[8][18]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[8][18]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[8][18]),
    .merge_data_o                                      (merge_data_pe_2_nw[8][18]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[8][18]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[8][18]),
    .gather_data_i                                     (gather_data_nw_2_pe[8][18]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[8][18]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[8][18]),
    .gather_data_o                                     (gather_data_pe_2_nw[8][18]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[8][18]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[8][18])
);


virtual_pe #(
    .cast_out                                          (cast_out_8_19),
    .merge_in                                          (merge_in_8_19),
    .merge_out                                         (merge_out_8_19),
    .gather_in                                         (gather_in_8_19),
    .gather_out                                        (gather_out_8_19),
    .x                                                 (8),
    .y                                                 (19)
)vpe_8_19(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[8][19]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[8][19]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[8][19]),
    .cast_data_o                                       (cast_data_pe_2_nw[8][19]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[8][19]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[8][19]),
    .merge_data_i                                      (merge_data_nw_2_pe[8][19]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[8][19]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[8][19]),
    .merge_data_o                                      (merge_data_pe_2_nw[8][19]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[8][19]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[8][19]),
    .gather_data_i                                     (gather_data_nw_2_pe[8][19]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[8][19]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[8][19]),
    .gather_data_o                                     (gather_data_pe_2_nw[8][19]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[8][19]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[8][19])
);


virtual_pe #(
    .cast_out                                          (cast_out_8_20),
    .merge_in                                          (merge_in_8_20),
    .merge_out                                         (merge_out_8_20),
    .gather_in                                         (gather_in_8_20),
    .gather_out                                        (gather_out_8_20),
    .x                                                 (8),
    .y                                                 (20)
)vpe_8_20(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[8][20]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[8][20]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[8][20]),
    .cast_data_o                                       (cast_data_pe_2_nw[8][20]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[8][20]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[8][20]),
    .merge_data_i                                      (merge_data_nw_2_pe[8][20]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[8][20]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[8][20]),
    .merge_data_o                                      (merge_data_pe_2_nw[8][20]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[8][20]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[8][20]),
    .gather_data_i                                     (gather_data_nw_2_pe[8][20]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[8][20]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[8][20]),
    .gather_data_o                                     (gather_data_pe_2_nw[8][20]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[8][20]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[8][20])
);


virtual_pe #(
    .cast_out                                          (cast_out_8_21),
    .merge_in                                          (merge_in_8_21),
    .merge_out                                         (merge_out_8_21),
    .gather_in                                         (gather_in_8_21),
    .gather_out                                        (gather_out_8_21),
    .x                                                 (8),
    .y                                                 (21)
)vpe_8_21(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[8][21]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[8][21]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[8][21]),
    .cast_data_o                                       (cast_data_pe_2_nw[8][21]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[8][21]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[8][21]),
    .merge_data_i                                      (merge_data_nw_2_pe[8][21]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[8][21]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[8][21]),
    .merge_data_o                                      (merge_data_pe_2_nw[8][21]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[8][21]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[8][21]),
    .gather_data_i                                     (gather_data_nw_2_pe[8][21]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[8][21]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[8][21]),
    .gather_data_o                                     (gather_data_pe_2_nw[8][21]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[8][21]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[8][21])
);


virtual_pe #(
    .cast_out                                          (cast_out_8_22),
    .merge_in                                          (merge_in_8_22),
    .merge_out                                         (merge_out_8_22),
    .gather_in                                         (gather_in_8_22),
    .gather_out                                        (gather_out_8_22),
    .x                                                 (8),
    .y                                                 (22)
)vpe_8_22(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[8][22]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[8][22]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[8][22]),
    .cast_data_o                                       (cast_data_pe_2_nw[8][22]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[8][22]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[8][22]),
    .merge_data_i                                      (merge_data_nw_2_pe[8][22]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[8][22]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[8][22]),
    .merge_data_o                                      (merge_data_pe_2_nw[8][22]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[8][22]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[8][22]),
    .gather_data_i                                     (gather_data_nw_2_pe[8][22]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[8][22]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[8][22]),
    .gather_data_o                                     (gather_data_pe_2_nw[8][22]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[8][22]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[8][22])
);


virtual_pe #(
    .cast_out                                          (cast_out_8_23),
    .merge_in                                          (merge_in_8_23),
    .merge_out                                         (merge_out_8_23),
    .gather_in                                         (gather_in_8_23),
    .gather_out                                        (gather_out_8_23),
    .x                                                 (8),
    .y                                                 (23)
)vpe_8_23(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[8][23]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[8][23]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[8][23]),
    .cast_data_o                                       (cast_data_pe_2_nw[8][23]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[8][23]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[8][23]),
    .merge_data_i                                      (merge_data_nw_2_pe[8][23]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[8][23]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[8][23]),
    .merge_data_o                                      (merge_data_pe_2_nw[8][23]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[8][23]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[8][23]),
    .gather_data_i                                     (gather_data_nw_2_pe[8][23]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[8][23]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[8][23]),
    .gather_data_o                                     (gather_data_pe_2_nw[8][23]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[8][23]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[8][23])
);


virtual_pe #(
    .cast_out                                          (cast_out_8_24),
    .merge_in                                          (merge_in_8_24),
    .merge_out                                         (merge_out_8_24),
    .gather_in                                         (gather_in_8_24),
    .gather_out                                        (gather_out_8_24),
    .x                                                 (8),
    .y                                                 (24)
)vpe_8_24(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[8][24]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[8][24]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[8][24]),
    .cast_data_o                                       (cast_data_pe_2_nw[8][24]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[8][24]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[8][24]),
    .merge_data_i                                      (merge_data_nw_2_pe[8][24]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[8][24]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[8][24]),
    .merge_data_o                                      (merge_data_pe_2_nw[8][24]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[8][24]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[8][24]),
    .gather_data_i                                     (gather_data_nw_2_pe[8][24]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[8][24]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[8][24]),
    .gather_data_o                                     (gather_data_pe_2_nw[8][24]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[8][24]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[8][24])
);


virtual_pe #(
    .cast_out                                          (cast_out_9_0),
    .merge_in                                          (merge_in_9_0),
    .merge_out                                         (merge_out_9_0),
    .gather_in                                         (gather_in_9_0),
    .gather_out                                        (gather_out_9_0),
    .x                                                 (9),
    .y                                                 (0)
)vpe_9_0(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[9][0]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[9][0]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[9][0]),
    .cast_data_o                                       (cast_data_pe_2_nw[9][0]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[9][0]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[9][0]),
    .merge_data_i                                      (merge_data_nw_2_pe[9][0]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[9][0]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[9][0]),
    .merge_data_o                                      (merge_data_pe_2_nw[9][0]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[9][0]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[9][0]),
    .gather_data_i                                     (gather_data_nw_2_pe[9][0]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[9][0]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[9][0]),
    .gather_data_o                                     (gather_data_pe_2_nw[9][0]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[9][0]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[9][0])
);


virtual_pe #(
    .cast_out                                          (cast_out_9_1),
    .merge_in                                          (merge_in_9_1),
    .merge_out                                         (merge_out_9_1),
    .gather_in                                         (gather_in_9_1),
    .gather_out                                        (gather_out_9_1),
    .x                                                 (9),
    .y                                                 (1)
)vpe_9_1(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[9][1]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[9][1]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[9][1]),
    .cast_data_o                                       (cast_data_pe_2_nw[9][1]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[9][1]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[9][1]),
    .merge_data_i                                      (merge_data_nw_2_pe[9][1]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[9][1]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[9][1]),
    .merge_data_o                                      (merge_data_pe_2_nw[9][1]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[9][1]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[9][1]),
    .gather_data_i                                     (gather_data_nw_2_pe[9][1]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[9][1]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[9][1]),
    .gather_data_o                                     (gather_data_pe_2_nw[9][1]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[9][1]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[9][1])
);


virtual_pe #(
    .cast_out                                          (cast_out_9_2),
    .merge_in                                          (merge_in_9_2),
    .merge_out                                         (merge_out_9_2),
    .gather_in                                         (gather_in_9_2),
    .gather_out                                        (gather_out_9_2),
    .x                                                 (9),
    .y                                                 (2)
)vpe_9_2(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[9][2]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[9][2]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[9][2]),
    .cast_data_o                                       (cast_data_pe_2_nw[9][2]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[9][2]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[9][2]),
    .merge_data_i                                      (merge_data_nw_2_pe[9][2]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[9][2]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[9][2]),
    .merge_data_o                                      (merge_data_pe_2_nw[9][2]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[9][2]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[9][2]),
    .gather_data_i                                     (gather_data_nw_2_pe[9][2]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[9][2]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[9][2]),
    .gather_data_o                                     (gather_data_pe_2_nw[9][2]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[9][2]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[9][2])
);


virtual_pe #(
    .cast_out                                          (cast_out_9_3),
    .merge_in                                          (merge_in_9_3),
    .merge_out                                         (merge_out_9_3),
    .gather_in                                         (gather_in_9_3),
    .gather_out                                        (gather_out_9_3),
    .x                                                 (9),
    .y                                                 (3)
)vpe_9_3(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[9][3]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[9][3]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[9][3]),
    .cast_data_o                                       (cast_data_pe_2_nw[9][3]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[9][3]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[9][3]),
    .merge_data_i                                      (merge_data_nw_2_pe[9][3]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[9][3]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[9][3]),
    .merge_data_o                                      (merge_data_pe_2_nw[9][3]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[9][3]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[9][3]),
    .gather_data_i                                     (gather_data_nw_2_pe[9][3]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[9][3]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[9][3]),
    .gather_data_o                                     (gather_data_pe_2_nw[9][3]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[9][3]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[9][3])
);


virtual_pe #(
    .cast_out                                          (cast_out_9_4),
    .merge_in                                          (merge_in_9_4),
    .merge_out                                         (merge_out_9_4),
    .gather_in                                         (gather_in_9_4),
    .gather_out                                        (gather_out_9_4),
    .x                                                 (9),
    .y                                                 (4)
)vpe_9_4(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[9][4]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[9][4]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[9][4]),
    .cast_data_o                                       (cast_data_pe_2_nw[9][4]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[9][4]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[9][4]),
    .merge_data_i                                      (merge_data_nw_2_pe[9][4]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[9][4]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[9][4]),
    .merge_data_o                                      (merge_data_pe_2_nw[9][4]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[9][4]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[9][4]),
    .gather_data_i                                     (gather_data_nw_2_pe[9][4]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[9][4]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[9][4]),
    .gather_data_o                                     (gather_data_pe_2_nw[9][4]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[9][4]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[9][4])
);


virtual_pe #(
    .cast_out                                          (cast_out_9_5),
    .merge_in                                          (merge_in_9_5),
    .merge_out                                         (merge_out_9_5),
    .gather_in                                         (gather_in_9_5),
    .gather_out                                        (gather_out_9_5),
    .x                                                 (9),
    .y                                                 (5)
)vpe_9_5(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[9][5]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[9][5]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[9][5]),
    .cast_data_o                                       (cast_data_pe_2_nw[9][5]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[9][5]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[9][5]),
    .merge_data_i                                      (merge_data_nw_2_pe[9][5]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[9][5]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[9][5]),
    .merge_data_o                                      (merge_data_pe_2_nw[9][5]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[9][5]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[9][5]),
    .gather_data_i                                     (gather_data_nw_2_pe[9][5]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[9][5]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[9][5]),
    .gather_data_o                                     (gather_data_pe_2_nw[9][5]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[9][5]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[9][5])
);


virtual_pe #(
    .cast_out                                          (cast_out_9_6),
    .merge_in                                          (merge_in_9_6),
    .merge_out                                         (merge_out_9_6),
    .gather_in                                         (gather_in_9_6),
    .gather_out                                        (gather_out_9_6),
    .x                                                 (9),
    .y                                                 (6)
)vpe_9_6(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[9][6]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[9][6]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[9][6]),
    .cast_data_o                                       (cast_data_pe_2_nw[9][6]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[9][6]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[9][6]),
    .merge_data_i                                      (merge_data_nw_2_pe[9][6]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[9][6]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[9][6]),
    .merge_data_o                                      (merge_data_pe_2_nw[9][6]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[9][6]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[9][6]),
    .gather_data_i                                     (gather_data_nw_2_pe[9][6]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[9][6]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[9][6]),
    .gather_data_o                                     (gather_data_pe_2_nw[9][6]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[9][6]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[9][6])
);


virtual_pe #(
    .cast_out                                          (cast_out_9_7),
    .merge_in                                          (merge_in_9_7),
    .merge_out                                         (merge_out_9_7),
    .gather_in                                         (gather_in_9_7),
    .gather_out                                        (gather_out_9_7),
    .x                                                 (9),
    .y                                                 (7)
)vpe_9_7(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[9][7]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[9][7]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[9][7]),
    .cast_data_o                                       (cast_data_pe_2_nw[9][7]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[9][7]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[9][7]),
    .merge_data_i                                      (merge_data_nw_2_pe[9][7]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[9][7]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[9][7]),
    .merge_data_o                                      (merge_data_pe_2_nw[9][7]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[9][7]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[9][7]),
    .gather_data_i                                     (gather_data_nw_2_pe[9][7]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[9][7]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[9][7]),
    .gather_data_o                                     (gather_data_pe_2_nw[9][7]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[9][7]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[9][7])
);


virtual_pe #(
    .cast_out                                          (cast_out_9_8),
    .merge_in                                          (merge_in_9_8),
    .merge_out                                         (merge_out_9_8),
    .gather_in                                         (gather_in_9_8),
    .gather_out                                        (gather_out_9_8),
    .x                                                 (9),
    .y                                                 (8)
)vpe_9_8(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[9][8]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[9][8]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[9][8]),
    .cast_data_o                                       (cast_data_pe_2_nw[9][8]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[9][8]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[9][8]),
    .merge_data_i                                      (merge_data_nw_2_pe[9][8]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[9][8]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[9][8]),
    .merge_data_o                                      (merge_data_pe_2_nw[9][8]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[9][8]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[9][8]),
    .gather_data_i                                     (gather_data_nw_2_pe[9][8]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[9][8]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[9][8]),
    .gather_data_o                                     (gather_data_pe_2_nw[9][8]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[9][8]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[9][8])
);


virtual_pe #(
    .cast_out                                          (cast_out_9_9),
    .merge_in                                          (merge_in_9_9),
    .merge_out                                         (merge_out_9_9),
    .gather_in                                         (gather_in_9_9),
    .gather_out                                        (gather_out_9_9),
    .x                                                 (9),
    .y                                                 (9)
)vpe_9_9(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[9][9]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[9][9]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[9][9]),
    .cast_data_o                                       (cast_data_pe_2_nw[9][9]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[9][9]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[9][9]),
    .merge_data_i                                      (merge_data_nw_2_pe[9][9]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[9][9]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[9][9]),
    .merge_data_o                                      (merge_data_pe_2_nw[9][9]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[9][9]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[9][9]),
    .gather_data_i                                     (gather_data_nw_2_pe[9][9]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[9][9]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[9][9]),
    .gather_data_o                                     (gather_data_pe_2_nw[9][9]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[9][9]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[9][9])
);


virtual_pe #(
    .cast_out                                          (cast_out_9_10),
    .merge_in                                          (merge_in_9_10),
    .merge_out                                         (merge_out_9_10),
    .gather_in                                         (gather_in_9_10),
    .gather_out                                        (gather_out_9_10),
    .x                                                 (9),
    .y                                                 (10)
)vpe_9_10(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[9][10]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[9][10]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[9][10]),
    .cast_data_o                                       (cast_data_pe_2_nw[9][10]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[9][10]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[9][10]),
    .merge_data_i                                      (merge_data_nw_2_pe[9][10]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[9][10]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[9][10]),
    .merge_data_o                                      (merge_data_pe_2_nw[9][10]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[9][10]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[9][10]),
    .gather_data_i                                     (gather_data_nw_2_pe[9][10]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[9][10]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[9][10]),
    .gather_data_o                                     (gather_data_pe_2_nw[9][10]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[9][10]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[9][10])
);


virtual_pe #(
    .cast_out                                          (cast_out_9_11),
    .merge_in                                          (merge_in_9_11),
    .merge_out                                         (merge_out_9_11),
    .gather_in                                         (gather_in_9_11),
    .gather_out                                        (gather_out_9_11),
    .x                                                 (9),
    .y                                                 (11)
)vpe_9_11(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[9][11]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[9][11]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[9][11]),
    .cast_data_o                                       (cast_data_pe_2_nw[9][11]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[9][11]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[9][11]),
    .merge_data_i                                      (merge_data_nw_2_pe[9][11]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[9][11]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[9][11]),
    .merge_data_o                                      (merge_data_pe_2_nw[9][11]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[9][11]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[9][11]),
    .gather_data_i                                     (gather_data_nw_2_pe[9][11]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[9][11]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[9][11]),
    .gather_data_o                                     (gather_data_pe_2_nw[9][11]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[9][11]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[9][11])
);


virtual_pe #(
    .cast_out                                          (cast_out_9_12),
    .merge_in                                          (merge_in_9_12),
    .merge_out                                         (merge_out_9_12),
    .gather_in                                         (gather_in_9_12),
    .gather_out                                        (gather_out_9_12),
    .x                                                 (9),
    .y                                                 (12)
)vpe_9_12(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[9][12]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[9][12]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[9][12]),
    .cast_data_o                                       (cast_data_pe_2_nw[9][12]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[9][12]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[9][12]),
    .merge_data_i                                      (merge_data_nw_2_pe[9][12]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[9][12]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[9][12]),
    .merge_data_o                                      (merge_data_pe_2_nw[9][12]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[9][12]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[9][12]),
    .gather_data_i                                     (gather_data_nw_2_pe[9][12]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[9][12]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[9][12]),
    .gather_data_o                                     (gather_data_pe_2_nw[9][12]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[9][12]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[9][12])
);


virtual_pe #(
    .cast_out                                          (cast_out_9_13),
    .merge_in                                          (merge_in_9_13),
    .merge_out                                         (merge_out_9_13),
    .gather_in                                         (gather_in_9_13),
    .gather_out                                        (gather_out_9_13),
    .x                                                 (9),
    .y                                                 (13)
)vpe_9_13(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[9][13]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[9][13]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[9][13]),
    .cast_data_o                                       (cast_data_pe_2_nw[9][13]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[9][13]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[9][13]),
    .merge_data_i                                      (merge_data_nw_2_pe[9][13]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[9][13]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[9][13]),
    .merge_data_o                                      (merge_data_pe_2_nw[9][13]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[9][13]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[9][13]),
    .gather_data_i                                     (gather_data_nw_2_pe[9][13]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[9][13]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[9][13]),
    .gather_data_o                                     (gather_data_pe_2_nw[9][13]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[9][13]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[9][13])
);


virtual_pe #(
    .cast_out                                          (cast_out_9_14),
    .merge_in                                          (merge_in_9_14),
    .merge_out                                         (merge_out_9_14),
    .gather_in                                         (gather_in_9_14),
    .gather_out                                        (gather_out_9_14),
    .x                                                 (9),
    .y                                                 (14)
)vpe_9_14(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[9][14]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[9][14]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[9][14]),
    .cast_data_o                                       (cast_data_pe_2_nw[9][14]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[9][14]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[9][14]),
    .merge_data_i                                      (merge_data_nw_2_pe[9][14]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[9][14]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[9][14]),
    .merge_data_o                                      (merge_data_pe_2_nw[9][14]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[9][14]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[9][14]),
    .gather_data_i                                     (gather_data_nw_2_pe[9][14]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[9][14]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[9][14]),
    .gather_data_o                                     (gather_data_pe_2_nw[9][14]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[9][14]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[9][14])
);


virtual_pe #(
    .cast_out                                          (cast_out_9_15),
    .merge_in                                          (merge_in_9_15),
    .merge_out                                         (merge_out_9_15),
    .gather_in                                         (gather_in_9_15),
    .gather_out                                        (gather_out_9_15),
    .x                                                 (9),
    .y                                                 (15)
)vpe_9_15(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[9][15]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[9][15]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[9][15]),
    .cast_data_o                                       (cast_data_pe_2_nw[9][15]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[9][15]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[9][15]),
    .merge_data_i                                      (merge_data_nw_2_pe[9][15]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[9][15]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[9][15]),
    .merge_data_o                                      (merge_data_pe_2_nw[9][15]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[9][15]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[9][15]),
    .gather_data_i                                     (gather_data_nw_2_pe[9][15]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[9][15]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[9][15]),
    .gather_data_o                                     (gather_data_pe_2_nw[9][15]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[9][15]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[9][15])
);


virtual_pe #(
    .cast_out                                          (cast_out_9_16),
    .merge_in                                          (merge_in_9_16),
    .merge_out                                         (merge_out_9_16),
    .gather_in                                         (gather_in_9_16),
    .gather_out                                        (gather_out_9_16),
    .x                                                 (9),
    .y                                                 (16)
)vpe_9_16(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[9][16]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[9][16]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[9][16]),
    .cast_data_o                                       (cast_data_pe_2_nw[9][16]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[9][16]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[9][16]),
    .merge_data_i                                      (merge_data_nw_2_pe[9][16]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[9][16]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[9][16]),
    .merge_data_o                                      (merge_data_pe_2_nw[9][16]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[9][16]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[9][16]),
    .gather_data_i                                     (gather_data_nw_2_pe[9][16]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[9][16]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[9][16]),
    .gather_data_o                                     (gather_data_pe_2_nw[9][16]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[9][16]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[9][16])
);


virtual_pe #(
    .cast_out                                          (cast_out_9_17),
    .merge_in                                          (merge_in_9_17),
    .merge_out                                         (merge_out_9_17),
    .gather_in                                         (gather_in_9_17),
    .gather_out                                        (gather_out_9_17),
    .x                                                 (9),
    .y                                                 (17)
)vpe_9_17(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[9][17]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[9][17]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[9][17]),
    .cast_data_o                                       (cast_data_pe_2_nw[9][17]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[9][17]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[9][17]),
    .merge_data_i                                      (merge_data_nw_2_pe[9][17]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[9][17]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[9][17]),
    .merge_data_o                                      (merge_data_pe_2_nw[9][17]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[9][17]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[9][17]),
    .gather_data_i                                     (gather_data_nw_2_pe[9][17]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[9][17]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[9][17]),
    .gather_data_o                                     (gather_data_pe_2_nw[9][17]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[9][17]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[9][17])
);


virtual_pe #(
    .cast_out                                          (cast_out_9_18),
    .merge_in                                          (merge_in_9_18),
    .merge_out                                         (merge_out_9_18),
    .gather_in                                         (gather_in_9_18),
    .gather_out                                        (gather_out_9_18),
    .x                                                 (9),
    .y                                                 (18)
)vpe_9_18(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[9][18]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[9][18]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[9][18]),
    .cast_data_o                                       (cast_data_pe_2_nw[9][18]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[9][18]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[9][18]),
    .merge_data_i                                      (merge_data_nw_2_pe[9][18]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[9][18]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[9][18]),
    .merge_data_o                                      (merge_data_pe_2_nw[9][18]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[9][18]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[9][18]),
    .gather_data_i                                     (gather_data_nw_2_pe[9][18]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[9][18]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[9][18]),
    .gather_data_o                                     (gather_data_pe_2_nw[9][18]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[9][18]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[9][18])
);


virtual_pe #(
    .cast_out                                          (cast_out_9_19),
    .merge_in                                          (merge_in_9_19),
    .merge_out                                         (merge_out_9_19),
    .gather_in                                         (gather_in_9_19),
    .gather_out                                        (gather_out_9_19),
    .x                                                 (9),
    .y                                                 (19)
)vpe_9_19(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[9][19]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[9][19]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[9][19]),
    .cast_data_o                                       (cast_data_pe_2_nw[9][19]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[9][19]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[9][19]),
    .merge_data_i                                      (merge_data_nw_2_pe[9][19]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[9][19]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[9][19]),
    .merge_data_o                                      (merge_data_pe_2_nw[9][19]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[9][19]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[9][19]),
    .gather_data_i                                     (gather_data_nw_2_pe[9][19]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[9][19]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[9][19]),
    .gather_data_o                                     (gather_data_pe_2_nw[9][19]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[9][19]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[9][19])
);


virtual_pe #(
    .cast_out                                          (cast_out_9_20),
    .merge_in                                          (merge_in_9_20),
    .merge_out                                         (merge_out_9_20),
    .gather_in                                         (gather_in_9_20),
    .gather_out                                        (gather_out_9_20),
    .x                                                 (9),
    .y                                                 (20)
)vpe_9_20(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[9][20]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[9][20]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[9][20]),
    .cast_data_o                                       (cast_data_pe_2_nw[9][20]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[9][20]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[9][20]),
    .merge_data_i                                      (merge_data_nw_2_pe[9][20]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[9][20]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[9][20]),
    .merge_data_o                                      (merge_data_pe_2_nw[9][20]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[9][20]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[9][20]),
    .gather_data_i                                     (gather_data_nw_2_pe[9][20]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[9][20]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[9][20]),
    .gather_data_o                                     (gather_data_pe_2_nw[9][20]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[9][20]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[9][20])
);


virtual_pe #(
    .cast_out                                          (cast_out_9_21),
    .merge_in                                          (merge_in_9_21),
    .merge_out                                         (merge_out_9_21),
    .gather_in                                         (gather_in_9_21),
    .gather_out                                        (gather_out_9_21),
    .x                                                 (9),
    .y                                                 (21)
)vpe_9_21(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[9][21]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[9][21]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[9][21]),
    .cast_data_o                                       (cast_data_pe_2_nw[9][21]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[9][21]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[9][21]),
    .merge_data_i                                      (merge_data_nw_2_pe[9][21]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[9][21]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[9][21]),
    .merge_data_o                                      (merge_data_pe_2_nw[9][21]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[9][21]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[9][21]),
    .gather_data_i                                     (gather_data_nw_2_pe[9][21]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[9][21]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[9][21]),
    .gather_data_o                                     (gather_data_pe_2_nw[9][21]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[9][21]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[9][21])
);


virtual_pe #(
    .cast_out                                          (cast_out_9_22),
    .merge_in                                          (merge_in_9_22),
    .merge_out                                         (merge_out_9_22),
    .gather_in                                         (gather_in_9_22),
    .gather_out                                        (gather_out_9_22),
    .x                                                 (9),
    .y                                                 (22)
)vpe_9_22(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[9][22]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[9][22]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[9][22]),
    .cast_data_o                                       (cast_data_pe_2_nw[9][22]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[9][22]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[9][22]),
    .merge_data_i                                      (merge_data_nw_2_pe[9][22]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[9][22]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[9][22]),
    .merge_data_o                                      (merge_data_pe_2_nw[9][22]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[9][22]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[9][22]),
    .gather_data_i                                     (gather_data_nw_2_pe[9][22]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[9][22]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[9][22]),
    .gather_data_o                                     (gather_data_pe_2_nw[9][22]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[9][22]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[9][22])
);


virtual_pe #(
    .cast_out                                          (cast_out_9_23),
    .merge_in                                          (merge_in_9_23),
    .merge_out                                         (merge_out_9_23),
    .gather_in                                         (gather_in_9_23),
    .gather_out                                        (gather_out_9_23),
    .x                                                 (9),
    .y                                                 (23)
)vpe_9_23(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[9][23]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[9][23]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[9][23]),
    .cast_data_o                                       (cast_data_pe_2_nw[9][23]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[9][23]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[9][23]),
    .merge_data_i                                      (merge_data_nw_2_pe[9][23]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[9][23]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[9][23]),
    .merge_data_o                                      (merge_data_pe_2_nw[9][23]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[9][23]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[9][23]),
    .gather_data_i                                     (gather_data_nw_2_pe[9][23]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[9][23]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[9][23]),
    .gather_data_o                                     (gather_data_pe_2_nw[9][23]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[9][23]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[9][23])
);


virtual_pe #(
    .cast_out                                          (cast_out_9_24),
    .merge_in                                          (merge_in_9_24),
    .merge_out                                         (merge_out_9_24),
    .gather_in                                         (gather_in_9_24),
    .gather_out                                        (gather_out_9_24),
    .x                                                 (9),
    .y                                                 (24)
)vpe_9_24(
    .clk                                               (clk),
    .rstn                                              (rstn),
    .cast_data_i                                       (cast_data_nw_2_pe[9][24]),
    .cast_valid_i                                      (cast_valid_nw_2_pe[9][24]),
    .cast_ready_o                                      (cast_ready_pe_2_nw[9][24]),
    .cast_data_o                                       (cast_data_pe_2_nw[9][24]),
    .cast_valid_o                                      (cast_valid_pe_2_nw[9][24]),
    .cast_ready_i                                      (cast_ready_nw_2_pe[9][24]),
    .merge_data_i                                      (merge_data_nw_2_pe[9][24]),
    .merge_valid_i                                     (merge_valid_nw_2_pe[9][24]),
    .merge_ready_o                                     (merge_ready_pe_2_nw[9][24]),
    .merge_data_o                                      (merge_data_pe_2_nw[9][24]),
    .merge_valid_o                                     (merge_valid_pe_2_nw[9][24]),
    .merge_ready_i                                     (merge_ready_nw_2_pe[9][24]),
    .gather_data_i                                     (gather_data_nw_2_pe[9][24]),
    .gather_valid_i                                    (gather_valid_nw_2_pe[9][24]),
    .gather_ready_o                                    (gather_ready_pe_2_nw[9][24]),
    .gather_data_o                                     (gather_data_pe_2_nw[9][24]),
    .gather_valid_o                                    (gather_valid_pe_2_nw[9][24]),
    .gather_ready_i                                    (gather_ready_nw_2_pe[9][24])
);

endmodule
