localparam isFC_list_0_0[`CN] = '{0,0,0,0,0};
localparam isFC_list_1_0[`CN] = '{0,0,0,0,0};
localparam isFC_list_2_0[`CN] = '{0,0,0,0,0};
localparam isFC_list_3_0[`CN] = '{0,0,0,0,0};
localparam isFC_list_4_0[`CN] = '{0,0,0,0,0};
localparam isFC_list_5_0[`CN] = '{0,0,0,0,0};
localparam isFC_list_6_0[`CN] = '{0,0,0,0,0};
localparam isFC_list_0_1[`CN] = '{0,0,0,0,0};
localparam isFC_list_1_1[`CN] = '{0,0,0,0,0};
localparam isFC_list_2_1[`CN] = '{0,0,0,0,0};
localparam isFC_list_3_1[`CN] = '{1,1,1,0,0};
localparam isFC_list_4_1[`CN] = '{0,0,0,0,0};
localparam isFC_list_5_1[`CN] = '{0,0,0,0,0};
localparam isFC_list_6_1[`CN] = '{0,0,0,0,0};
localparam isFC_list_0_2[`CN] = '{0,0,0,0,0};
localparam isFC_list_1_2[`CN] = '{0,0,0,0,0};
localparam isFC_list_2_2[`CN] = '{0,0,0,0,0};
localparam isFC_list_3_2[`CN] = '{0,0,0,0,0};
localparam isFC_list_4_2[`CN] = '{0,0,0,0,0};
localparam isFC_list_5_2[`CN] = '{0,0,0,0,0};
localparam isFC_list_6_2[`CN] = '{0,0,0,0,0};
localparam isFC_list_1_3[`CN] = '{0,0,0,0,0};
localparam isFC_list_0_3[`CN] = '{0,0,0,0,0};
localparam isFC_list_1_3[`CN] = '{0,0,0,0,0};
localparam isFC_list_2_3[`CN] = '{0,0,0,0,0};
localparam isFC_list_3_3[`CN] = '{0,0,0,0,0};
localparam isFC_list_4_3[`CN] = '{0,0,0,0,0};
localparam isFC_list_5_3[`CN] = '{0,0,0,0,0};
localparam isFC_list_6_4[`CN] = '{0,0,0,0,0};
localparam isFC_list_1_4[`CN] = '{0,0,0,0,0};
localparam isFC_list_2_4[`CN] = '{1,1,0,0,0};
localparam isFC_list_3_4[`CN] = '{0,0,0,0,0};
localparam isFC_list_4_4[`CN] = '{0,0,0,0,0};
localparam isFC_list_5_4[`CN] = '{0,0,0,0,0};
localparam isFC_list_6_4[`CN] = '{0,0,0,0,0};
localparam isFC_list_0_5[`CN] = '{0,0,0,0,0};
localparam isFC_list_1_5[`CN] = '{0,0,0,0,0};
localparam isFC_list_2_5[`CN] = '{0,0,0,0,0};
localparam isFC_list_3_5[`CN] = '{0,0,0,0,0};
localparam isFC_list_4_5[`CN] = '{0,0,0,0,0};
localparam isFC_list_5_5[`CN] = '{0,0,0,0,0};
localparam isFC_list_6_5[`CN] = '{0,0,0,0,0};
localparam isFC_list_0_6[`CN] = '{0,0,0,0,0};
localparam isFC_list_1_6[`CN] = '{0,0,0,0,0};
localparam isFC_list_2_6[`CN] = '{0,0,0,0,0};
localparam isFC_list_3_6[`CN] = '{0,0,0,0,0};
localparam isFC_list_4_6[`CN] = '{0,0,0,0,0};
localparam isFC_list_5_6[`CN] = '{0,0,0,0,0};
localparam isFC_list_6_6[`CN] = '{0,0,0,0,0};
localparam isFC_list_0_7[`CN] = '{0,0,0,0,0};
localparam isFC_list_1_7[`CN] = '{0,0,0,0,0};
localparam isFC_list_2_7[`CN] = '{1,1,0,0,0};
localparam isFC_list_3_7[`CN] = '{0,0,0,0,0};
localparam isFC_list_4_7[`CN] = '{0,0,0,0,0};
localparam isFC_list_5_7[`CN] = '{0,0,0,0,0};
localparam isFC_list_6_7[`CN] = '{0,0,0,0,0};

localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_0_0[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_1_0[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_2_0[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};//note the reverse index
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_3_0[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_4_0[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_5_0[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_6_0[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_0_1[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_1_1[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_2_1[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_3_1[`CN] = '{56'b00000000000000000000000000000000000110011000000000000000,56'b00000000000000000000000000000000000001100000000000000000,56'b00000000000000000000000000000000000000000000011100000000,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_4_1[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_5_1[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_6_1[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_0_2[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_1_2[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_2_2[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_3_2[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_4_2[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_5_2[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_6_2[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_0_3[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_1_3[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_2_3[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_3_3[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_4_3[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_5_3[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_6_3[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_0_4[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_1_4[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_2_4[`CN] = '{56'b00000000000000001101100000000000000000000000000000000000,56'b00000000000000110000000110000000000000000000000000000000,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_3_4[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_4_4[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_5_4[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_6_4[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_0_5[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_1_5[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_2_5[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_3_5[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_4_5[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_5_5[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_6_5[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_0_6[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_1_6[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_2_6[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_3_6[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_4_6[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_5_6[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_6_6[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_0_7[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_1_7[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_2_7[`CN] = '{56'b11110000000000000000000000000000000000000000000000000000,56'b00000001111000000000000000000000000000000000000000000000,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_3_7[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_4_7[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_5_7[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_6_7[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};

localparam int FCpl_list_0_0[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_1_0[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_2_0[`CN] = '{16,0,0,0,0};
localparam int FCpl_list_0_1[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_1_1[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_2_1[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_0_2[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_1_2[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_2_2[`CN] = '{0,0,0,0,0};

localparam string rt_file_list_0_0[`CN] = '{"/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_0_0_0","/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_0_0_1","/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_0_0_2","/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_0_0_3","/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_0_0_4"};
localparam string rt_file_list_1_0[`CN] = '{"/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_1_0_0","/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_1_0_1","/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_1_0_2","/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_1_0_3","/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_1_0_4"};
localparam string rt_file_list_2_0[`CN] = '{"/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_2_0_0","/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_2_0_1","/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_2_0_2","/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_2_0_3","/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_2_0_4"};
localparam string rt_file_list_0_1[`CN] = '{"/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_0_1_0","/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_0_1_1","/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_0_1_2","/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_0_1_3","/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_0_1_4"};
localparam string rt_file_list_1_1[`CN] = '{"/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_1_1_0","/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_1_1_1","/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_1_1_2","/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_1_1_3","/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_1_1_4"};
localparam string rt_file_list_2_1[`CN] = '{"/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_2_1_0","/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_2_1_1","/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_2_1_2","/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_2_1_3","/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_2_1_4"};
localparam string rt_file_list_0_2[`CN] = '{"/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_0_2_0","/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_0_2_1","/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_0_2_2","/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_0_2_3","/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_0_2_4"};
localparam string rt_file_list_1_2[`CN] = '{"/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_1_2_0","/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_1_2_1","/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_1_2_2","/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_1_2_3","/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_1_2_4"};
localparam string rt_file_list_2_2[`CN] = '{"/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_2_2_0","/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_2_2_1","/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_2_2_2","/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_2_2_3","/mnt/c/git/NVCIM-COMM/behavior_model/test_multicast/config/cast_rt_2_2_4"};
