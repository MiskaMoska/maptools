`include "params.svh"
`include "network_config.svh"

module network(
    input       wire                        clk,
    input       wire                        rstn,

    //stab port
    input       wire        [`DW-1:0]       data_i_stab,
    input       wire                        valid_i_stab,
    output      wire                        ready_o_stab,

    //flee0 port
    output      wire        [`DW-1:0]       data_o_flee0,
    output      wire                        valid_o_flee0,
    input       wire                        ready_i_flee0,

    //flee1 port
    output      wire        [`DW-1:0]       data_o_flee1,
    output      wire                        valid_o_flee1,
    input       wire                        ready_i_flee1,

    //flee2 port
    output      wire        [`DW-1:0]       data_o_flee2,
    output      wire                        valid_o_flee2,
    input       wire                        ready_i_flee2,

    //flee3 port
    output      wire        [`DW-1:0]       data_o_flee3,
    output      wire                        valid_o_flee3,
    input       wire                        ready_i_flee3,

    //flee4 port
    output      wire        [`DW-1:0]       data_o_flee4,
    output      wire                        valid_o_flee4,
    input       wire                        ready_i_flee4,

    //flee5 port
    output      wire        [`DW-1:0]       data_o_flee5,
    output      wire                        valid_o_flee5,
    input       wire                        ready_i_flee5,

    //flee6 port
    output      wire        [`DW-1:0]       data_o_flee6,
    output      wire                        valid_o_flee6,
    input       wire                        ready_i_flee6,

    //flee7 port
    output      wire        [`DW-1:0]       data_o_flee7,
    output      wire                        valid_o_flee7,
    input       wire                        ready_i_flee7,

    input       wire        [`DW-1:0]       cast_data_i_0_0,
    input       wire                        cast_valid_i_0_0,
    output      wire                        cast_ready_o_0_0,

    output      wire        [`DW-1:0]       cast_data_o_0_0,
    output      wire                        cast_valid_o_0_0,
    input       wire                        cast_ready_i_0_0,

    input       wire        [`DW-1:0]       cast_data_i_0_1,
    input       wire                        cast_valid_i_0_1,
    output      wire                        cast_ready_o_0_1,

    output      wire        [`DW-1:0]       cast_data_o_0_1,
    output      wire                        cast_valid_o_0_1,
    input       wire                        cast_ready_i_0_1,

    input       wire        [`DW-1:0]       cast_data_i_0_2,
    input       wire                        cast_valid_i_0_2,
    output      wire                        cast_ready_o_0_2,

    output      wire        [`DW-1:0]       cast_data_o_0_2,
    output      wire                        cast_valid_o_0_2,
    input       wire                        cast_ready_i_0_2,

    input       wire        [`DW-1:0]       cast_data_i_0_3,
    input       wire                        cast_valid_i_0_3,
    output      wire                        cast_ready_o_0_3,

    output      wire        [`DW-1:0]       cast_data_o_0_3,
    output      wire                        cast_valid_o_0_3,
    input       wire                        cast_ready_i_0_3,

    input       wire        [`DW-1:0]       cast_data_i_0_4,
    input       wire                        cast_valid_i_0_4,
    output      wire                        cast_ready_o_0_4,

    output      wire        [`DW-1:0]       cast_data_o_0_4,
    output      wire                        cast_valid_o_0_4,
    input       wire                        cast_ready_i_0_4,

    input       wire        [`DW-1:0]       cast_data_i_0_5,
    input       wire                        cast_valid_i_0_5,
    output      wire                        cast_ready_o_0_5,

    output      wire        [`DW-1:0]       cast_data_o_0_5,
    output      wire                        cast_valid_o_0_5,
    input       wire                        cast_ready_i_0_5,

    input       wire        [`DW-1:0]       cast_data_i_0_6,
    input       wire                        cast_valid_i_0_6,
    output      wire                        cast_ready_o_0_6,

    output      wire        [`DW-1:0]       cast_data_o_0_6,
    output      wire                        cast_valid_o_0_6,
    input       wire                        cast_ready_i_0_6,

    input       wire        [`DW-1:0]       cast_data_i_0_7,
    input       wire                        cast_valid_i_0_7,
    output      wire                        cast_ready_o_0_7,

    output      wire        [`DW-1:0]       cast_data_o_0_7,
    output      wire                        cast_valid_o_0_7,
    input       wire                        cast_ready_i_0_7,

    input       wire        [`DW-1:0]       cast_data_i_0_8,
    input       wire                        cast_valid_i_0_8,
    output      wire                        cast_ready_o_0_8,

    output      wire        [`DW-1:0]       cast_data_o_0_8,
    output      wire                        cast_valid_o_0_8,
    input       wire                        cast_ready_i_0_8,

    input       wire        [`DW-1:0]       cast_data_i_0_9,
    input       wire                        cast_valid_i_0_9,
    output      wire                        cast_ready_o_0_9,

    output      wire        [`DW-1:0]       cast_data_o_0_9,
    output      wire                        cast_valid_o_0_9,
    input       wire                        cast_ready_i_0_9,

    input       wire        [`DW-1:0]       cast_data_i_0_10,
    input       wire                        cast_valid_i_0_10,
    output      wire                        cast_ready_o_0_10,

    output      wire        [`DW-1:0]       cast_data_o_0_10,
    output      wire                        cast_valid_o_0_10,
    input       wire                        cast_ready_i_0_10,

    input       wire        [`DW-1:0]       cast_data_i_0_11,
    input       wire                        cast_valid_i_0_11,
    output      wire                        cast_ready_o_0_11,

    output      wire        [`DW-1:0]       cast_data_o_0_11,
    output      wire                        cast_valid_o_0_11,
    input       wire                        cast_ready_i_0_11,

    input       wire        [`DW-1:0]       cast_data_i_0_12,
    input       wire                        cast_valid_i_0_12,
    output      wire                        cast_ready_o_0_12,

    output      wire        [`DW-1:0]       cast_data_o_0_12,
    output      wire                        cast_valid_o_0_12,
    input       wire                        cast_ready_i_0_12,

    input       wire        [`DW-1:0]       cast_data_i_0_13,
    input       wire                        cast_valid_i_0_13,
    output      wire                        cast_ready_o_0_13,

    output      wire        [`DW-1:0]       cast_data_o_0_13,
    output      wire                        cast_valid_o_0_13,
    input       wire                        cast_ready_i_0_13,

    input       wire        [`DW-1:0]       cast_data_i_0_14,
    input       wire                        cast_valid_i_0_14,
    output      wire                        cast_ready_o_0_14,

    output      wire        [`DW-1:0]       cast_data_o_0_14,
    output      wire                        cast_valid_o_0_14,
    input       wire                        cast_ready_i_0_14,

    input       wire        [`DW-1:0]       cast_data_i_0_15,
    input       wire                        cast_valid_i_0_15,
    output      wire                        cast_ready_o_0_15,

    output      wire        [`DW-1:0]       cast_data_o_0_15,
    output      wire                        cast_valid_o_0_15,
    input       wire                        cast_ready_i_0_15,

    input       wire        [`DW-1:0]       cast_data_i_0_16,
    input       wire                        cast_valid_i_0_16,
    output      wire                        cast_ready_o_0_16,

    output      wire        [`DW-1:0]       cast_data_o_0_16,
    output      wire                        cast_valid_o_0_16,
    input       wire                        cast_ready_i_0_16,

    input       wire        [`DW-1:0]       cast_data_i_0_17,
    input       wire                        cast_valid_i_0_17,
    output      wire                        cast_ready_o_0_17,

    output      wire        [`DW-1:0]       cast_data_o_0_17,
    output      wire                        cast_valid_o_0_17,
    input       wire                        cast_ready_i_0_17,

    input       wire        [`DW-1:0]       cast_data_i_0_18,
    input       wire                        cast_valid_i_0_18,
    output      wire                        cast_ready_o_0_18,

    output      wire        [`DW-1:0]       cast_data_o_0_18,
    output      wire                        cast_valid_o_0_18,
    input       wire                        cast_ready_i_0_18,

    input       wire        [`DW-1:0]       cast_data_i_0_19,
    input       wire                        cast_valid_i_0_19,
    output      wire                        cast_ready_o_0_19,

    output      wire        [`DW-1:0]       cast_data_o_0_19,
    output      wire                        cast_valid_o_0_19,
    input       wire                        cast_ready_i_0_19,

    input       wire        [`DW-1:0]       cast_data_i_0_20,
    input       wire                        cast_valid_i_0_20,
    output      wire                        cast_ready_o_0_20,

    output      wire        [`DW-1:0]       cast_data_o_0_20,
    output      wire                        cast_valid_o_0_20,
    input       wire                        cast_ready_i_0_20,

    input       wire        [`DW-1:0]       cast_data_i_0_21,
    input       wire                        cast_valid_i_0_21,
    output      wire                        cast_ready_o_0_21,

    output      wire        [`DW-1:0]       cast_data_o_0_21,
    output      wire                        cast_valid_o_0_21,
    input       wire                        cast_ready_i_0_21,

    input       wire        [`DW-1:0]       cast_data_i_0_22,
    input       wire                        cast_valid_i_0_22,
    output      wire                        cast_ready_o_0_22,

    output      wire        [`DW-1:0]       cast_data_o_0_22,
    output      wire                        cast_valid_o_0_22,
    input       wire                        cast_ready_i_0_22,

    input       wire        [`DW-1:0]       cast_data_i_0_23,
    input       wire                        cast_valid_i_0_23,
    output      wire                        cast_ready_o_0_23,

    output      wire        [`DW-1:0]       cast_data_o_0_23,
    output      wire                        cast_valid_o_0_23,
    input       wire                        cast_ready_i_0_23,

    input       wire        [`DW-1:0]       cast_data_i_0_24,
    input       wire                        cast_valid_i_0_24,
    output      wire                        cast_ready_o_0_24,

    output      wire        [`DW-1:0]       cast_data_o_0_24,
    output      wire                        cast_valid_o_0_24,
    input       wire                        cast_ready_i_0_24,

    input       wire        [`DW-1:0]       cast_data_i_1_0,
    input       wire                        cast_valid_i_1_0,
    output      wire                        cast_ready_o_1_0,

    output      wire        [`DW-1:0]       cast_data_o_1_0,
    output      wire                        cast_valid_o_1_0,
    input       wire                        cast_ready_i_1_0,

    input       wire        [`DW-1:0]       cast_data_i_1_1,
    input       wire                        cast_valid_i_1_1,
    output      wire                        cast_ready_o_1_1,

    output      wire        [`DW-1:0]       cast_data_o_1_1,
    output      wire                        cast_valid_o_1_1,
    input       wire                        cast_ready_i_1_1,

    input       wire        [`DW-1:0]       cast_data_i_1_2,
    input       wire                        cast_valid_i_1_2,
    output      wire                        cast_ready_o_1_2,

    output      wire        [`DW-1:0]       cast_data_o_1_2,
    output      wire                        cast_valid_o_1_2,
    input       wire                        cast_ready_i_1_2,

    input       wire        [`DW-1:0]       cast_data_i_1_3,
    input       wire                        cast_valid_i_1_3,
    output      wire                        cast_ready_o_1_3,

    output      wire        [`DW-1:0]       cast_data_o_1_3,
    output      wire                        cast_valid_o_1_3,
    input       wire                        cast_ready_i_1_3,

    input       wire        [`DW-1:0]       cast_data_i_1_4,
    input       wire                        cast_valid_i_1_4,
    output      wire                        cast_ready_o_1_4,

    output      wire        [`DW-1:0]       cast_data_o_1_4,
    output      wire                        cast_valid_o_1_4,
    input       wire                        cast_ready_i_1_4,

    input       wire        [`DW-1:0]       cast_data_i_1_5,
    input       wire                        cast_valid_i_1_5,
    output      wire                        cast_ready_o_1_5,

    output      wire        [`DW-1:0]       cast_data_o_1_5,
    output      wire                        cast_valid_o_1_5,
    input       wire                        cast_ready_i_1_5,

    input       wire        [`DW-1:0]       cast_data_i_1_6,
    input       wire                        cast_valid_i_1_6,
    output      wire                        cast_ready_o_1_6,

    output      wire        [`DW-1:0]       cast_data_o_1_6,
    output      wire                        cast_valid_o_1_6,
    input       wire                        cast_ready_i_1_6,

    input       wire        [`DW-1:0]       cast_data_i_1_7,
    input       wire                        cast_valid_i_1_7,
    output      wire                        cast_ready_o_1_7,

    output      wire        [`DW-1:0]       cast_data_o_1_7,
    output      wire                        cast_valid_o_1_7,
    input       wire                        cast_ready_i_1_7,

    input       wire        [`DW-1:0]       cast_data_i_1_8,
    input       wire                        cast_valid_i_1_8,
    output      wire                        cast_ready_o_1_8,

    output      wire        [`DW-1:0]       cast_data_o_1_8,
    output      wire                        cast_valid_o_1_8,
    input       wire                        cast_ready_i_1_8,

    input       wire        [`DW-1:0]       cast_data_i_1_9,
    input       wire                        cast_valid_i_1_9,
    output      wire                        cast_ready_o_1_9,

    output      wire        [`DW-1:0]       cast_data_o_1_9,
    output      wire                        cast_valid_o_1_9,
    input       wire                        cast_ready_i_1_9,

    input       wire        [`DW-1:0]       cast_data_i_1_10,
    input       wire                        cast_valid_i_1_10,
    output      wire                        cast_ready_o_1_10,

    output      wire        [`DW-1:0]       cast_data_o_1_10,
    output      wire                        cast_valid_o_1_10,
    input       wire                        cast_ready_i_1_10,

    input       wire        [`DW-1:0]       cast_data_i_1_11,
    input       wire                        cast_valid_i_1_11,
    output      wire                        cast_ready_o_1_11,

    output      wire        [`DW-1:0]       cast_data_o_1_11,
    output      wire                        cast_valid_o_1_11,
    input       wire                        cast_ready_i_1_11,

    input       wire        [`DW-1:0]       cast_data_i_1_12,
    input       wire                        cast_valid_i_1_12,
    output      wire                        cast_ready_o_1_12,

    output      wire        [`DW-1:0]       cast_data_o_1_12,
    output      wire                        cast_valid_o_1_12,
    input       wire                        cast_ready_i_1_12,

    input       wire        [`DW-1:0]       cast_data_i_1_13,
    input       wire                        cast_valid_i_1_13,
    output      wire                        cast_ready_o_1_13,

    output      wire        [`DW-1:0]       cast_data_o_1_13,
    output      wire                        cast_valid_o_1_13,
    input       wire                        cast_ready_i_1_13,

    input       wire        [`DW-1:0]       cast_data_i_1_14,
    input       wire                        cast_valid_i_1_14,
    output      wire                        cast_ready_o_1_14,

    output      wire        [`DW-1:0]       cast_data_o_1_14,
    output      wire                        cast_valid_o_1_14,
    input       wire                        cast_ready_i_1_14,

    input       wire        [`DW-1:0]       cast_data_i_1_15,
    input       wire                        cast_valid_i_1_15,
    output      wire                        cast_ready_o_1_15,

    output      wire        [`DW-1:0]       cast_data_o_1_15,
    output      wire                        cast_valid_o_1_15,
    input       wire                        cast_ready_i_1_15,

    input       wire        [`DW-1:0]       cast_data_i_1_16,
    input       wire                        cast_valid_i_1_16,
    output      wire                        cast_ready_o_1_16,

    output      wire        [`DW-1:0]       cast_data_o_1_16,
    output      wire                        cast_valid_o_1_16,
    input       wire                        cast_ready_i_1_16,

    input       wire        [`DW-1:0]       cast_data_i_1_17,
    input       wire                        cast_valid_i_1_17,
    output      wire                        cast_ready_o_1_17,

    output      wire        [`DW-1:0]       cast_data_o_1_17,
    output      wire                        cast_valid_o_1_17,
    input       wire                        cast_ready_i_1_17,

    input       wire        [`DW-1:0]       cast_data_i_1_18,
    input       wire                        cast_valid_i_1_18,
    output      wire                        cast_ready_o_1_18,

    output      wire        [`DW-1:0]       cast_data_o_1_18,
    output      wire                        cast_valid_o_1_18,
    input       wire                        cast_ready_i_1_18,

    input       wire        [`DW-1:0]       cast_data_i_1_19,
    input       wire                        cast_valid_i_1_19,
    output      wire                        cast_ready_o_1_19,

    output      wire        [`DW-1:0]       cast_data_o_1_19,
    output      wire                        cast_valid_o_1_19,
    input       wire                        cast_ready_i_1_19,

    input       wire        [`DW-1:0]       cast_data_i_1_20,
    input       wire                        cast_valid_i_1_20,
    output      wire                        cast_ready_o_1_20,

    output      wire        [`DW-1:0]       cast_data_o_1_20,
    output      wire                        cast_valid_o_1_20,
    input       wire                        cast_ready_i_1_20,

    input       wire        [`DW-1:0]       cast_data_i_1_21,
    input       wire                        cast_valid_i_1_21,
    output      wire                        cast_ready_o_1_21,

    output      wire        [`DW-1:0]       cast_data_o_1_21,
    output      wire                        cast_valid_o_1_21,
    input       wire                        cast_ready_i_1_21,

    input       wire        [`DW-1:0]       cast_data_i_1_22,
    input       wire                        cast_valid_i_1_22,
    output      wire                        cast_ready_o_1_22,

    output      wire        [`DW-1:0]       cast_data_o_1_22,
    output      wire                        cast_valid_o_1_22,
    input       wire                        cast_ready_i_1_22,

    input       wire        [`DW-1:0]       cast_data_i_1_23,
    input       wire                        cast_valid_i_1_23,
    output      wire                        cast_ready_o_1_23,

    output      wire        [`DW-1:0]       cast_data_o_1_23,
    output      wire                        cast_valid_o_1_23,
    input       wire                        cast_ready_i_1_23,

    input       wire        [`DW-1:0]       cast_data_i_1_24,
    input       wire                        cast_valid_i_1_24,
    output      wire                        cast_ready_o_1_24,

    output      wire        [`DW-1:0]       cast_data_o_1_24,
    output      wire                        cast_valid_o_1_24,
    input       wire                        cast_ready_i_1_24,

    input       wire        [`DW-1:0]       cast_data_i_2_0,
    input       wire                        cast_valid_i_2_0,
    output      wire                        cast_ready_o_2_0,

    output      wire        [`DW-1:0]       cast_data_o_2_0,
    output      wire                        cast_valid_o_2_0,
    input       wire                        cast_ready_i_2_0,

    input       wire        [`DW-1:0]       cast_data_i_2_1,
    input       wire                        cast_valid_i_2_1,
    output      wire                        cast_ready_o_2_1,

    output      wire        [`DW-1:0]       cast_data_o_2_1,
    output      wire                        cast_valid_o_2_1,
    input       wire                        cast_ready_i_2_1,

    input       wire        [`DW-1:0]       cast_data_i_2_2,
    input       wire                        cast_valid_i_2_2,
    output      wire                        cast_ready_o_2_2,

    output      wire        [`DW-1:0]       cast_data_o_2_2,
    output      wire                        cast_valid_o_2_2,
    input       wire                        cast_ready_i_2_2,

    input       wire        [`DW-1:0]       cast_data_i_2_3,
    input       wire                        cast_valid_i_2_3,
    output      wire                        cast_ready_o_2_3,

    output      wire        [`DW-1:0]       cast_data_o_2_3,
    output      wire                        cast_valid_o_2_3,
    input       wire                        cast_ready_i_2_3,

    input       wire        [`DW-1:0]       cast_data_i_2_4,
    input       wire                        cast_valid_i_2_4,
    output      wire                        cast_ready_o_2_4,

    output      wire        [`DW-1:0]       cast_data_o_2_4,
    output      wire                        cast_valid_o_2_4,
    input       wire                        cast_ready_i_2_4,

    input       wire        [`DW-1:0]       cast_data_i_2_5,
    input       wire                        cast_valid_i_2_5,
    output      wire                        cast_ready_o_2_5,

    output      wire        [`DW-1:0]       cast_data_o_2_5,
    output      wire                        cast_valid_o_2_5,
    input       wire                        cast_ready_i_2_5,

    input       wire        [`DW-1:0]       cast_data_i_2_6,
    input       wire                        cast_valid_i_2_6,
    output      wire                        cast_ready_o_2_6,

    output      wire        [`DW-1:0]       cast_data_o_2_6,
    output      wire                        cast_valid_o_2_6,
    input       wire                        cast_ready_i_2_6,

    input       wire        [`DW-1:0]       cast_data_i_2_7,
    input       wire                        cast_valid_i_2_7,
    output      wire                        cast_ready_o_2_7,

    output      wire        [`DW-1:0]       cast_data_o_2_7,
    output      wire                        cast_valid_o_2_7,
    input       wire                        cast_ready_i_2_7,

    input       wire        [`DW-1:0]       cast_data_i_2_8,
    input       wire                        cast_valid_i_2_8,
    output      wire                        cast_ready_o_2_8,

    output      wire        [`DW-1:0]       cast_data_o_2_8,
    output      wire                        cast_valid_o_2_8,
    input       wire                        cast_ready_i_2_8,

    input       wire        [`DW-1:0]       cast_data_i_2_9,
    input       wire                        cast_valid_i_2_9,
    output      wire                        cast_ready_o_2_9,

    output      wire        [`DW-1:0]       cast_data_o_2_9,
    output      wire                        cast_valid_o_2_9,
    input       wire                        cast_ready_i_2_9,

    input       wire        [`DW-1:0]       cast_data_i_2_10,
    input       wire                        cast_valid_i_2_10,
    output      wire                        cast_ready_o_2_10,

    output      wire        [`DW-1:0]       cast_data_o_2_10,
    output      wire                        cast_valid_o_2_10,
    input       wire                        cast_ready_i_2_10,

    input       wire        [`DW-1:0]       cast_data_i_2_11,
    input       wire                        cast_valid_i_2_11,
    output      wire                        cast_ready_o_2_11,

    output      wire        [`DW-1:0]       cast_data_o_2_11,
    output      wire                        cast_valid_o_2_11,
    input       wire                        cast_ready_i_2_11,

    input       wire        [`DW-1:0]       cast_data_i_2_12,
    input       wire                        cast_valid_i_2_12,
    output      wire                        cast_ready_o_2_12,

    output      wire        [`DW-1:0]       cast_data_o_2_12,
    output      wire                        cast_valid_o_2_12,
    input       wire                        cast_ready_i_2_12,

    input       wire        [`DW-1:0]       cast_data_i_2_13,
    input       wire                        cast_valid_i_2_13,
    output      wire                        cast_ready_o_2_13,

    output      wire        [`DW-1:0]       cast_data_o_2_13,
    output      wire                        cast_valid_o_2_13,
    input       wire                        cast_ready_i_2_13,

    input       wire        [`DW-1:0]       cast_data_i_2_14,
    input       wire                        cast_valid_i_2_14,
    output      wire                        cast_ready_o_2_14,

    output      wire        [`DW-1:0]       cast_data_o_2_14,
    output      wire                        cast_valid_o_2_14,
    input       wire                        cast_ready_i_2_14,

    input       wire        [`DW-1:0]       cast_data_i_2_15,
    input       wire                        cast_valid_i_2_15,
    output      wire                        cast_ready_o_2_15,

    output      wire        [`DW-1:0]       cast_data_o_2_15,
    output      wire                        cast_valid_o_2_15,
    input       wire                        cast_ready_i_2_15,

    input       wire        [`DW-1:0]       cast_data_i_2_16,
    input       wire                        cast_valid_i_2_16,
    output      wire                        cast_ready_o_2_16,

    output      wire        [`DW-1:0]       cast_data_o_2_16,
    output      wire                        cast_valid_o_2_16,
    input       wire                        cast_ready_i_2_16,

    input       wire        [`DW-1:0]       cast_data_i_2_17,
    input       wire                        cast_valid_i_2_17,
    output      wire                        cast_ready_o_2_17,

    output      wire        [`DW-1:0]       cast_data_o_2_17,
    output      wire                        cast_valid_o_2_17,
    input       wire                        cast_ready_i_2_17,

    input       wire        [`DW-1:0]       cast_data_i_2_18,
    input       wire                        cast_valid_i_2_18,
    output      wire                        cast_ready_o_2_18,

    output      wire        [`DW-1:0]       cast_data_o_2_18,
    output      wire                        cast_valid_o_2_18,
    input       wire                        cast_ready_i_2_18,

    input       wire        [`DW-1:0]       cast_data_i_2_19,
    input       wire                        cast_valid_i_2_19,
    output      wire                        cast_ready_o_2_19,

    output      wire        [`DW-1:0]       cast_data_o_2_19,
    output      wire                        cast_valid_o_2_19,
    input       wire                        cast_ready_i_2_19,

    input       wire        [`DW-1:0]       cast_data_i_2_20,
    input       wire                        cast_valid_i_2_20,
    output      wire                        cast_ready_o_2_20,

    output      wire        [`DW-1:0]       cast_data_o_2_20,
    output      wire                        cast_valid_o_2_20,
    input       wire                        cast_ready_i_2_20,

    input       wire        [`DW-1:0]       cast_data_i_2_21,
    input       wire                        cast_valid_i_2_21,
    output      wire                        cast_ready_o_2_21,

    output      wire        [`DW-1:0]       cast_data_o_2_21,
    output      wire                        cast_valid_o_2_21,
    input       wire                        cast_ready_i_2_21,

    input       wire        [`DW-1:0]       cast_data_i_2_22,
    input       wire                        cast_valid_i_2_22,
    output      wire                        cast_ready_o_2_22,

    output      wire        [`DW-1:0]       cast_data_o_2_22,
    output      wire                        cast_valid_o_2_22,
    input       wire                        cast_ready_i_2_22,

    input       wire        [`DW-1:0]       cast_data_i_2_23,
    input       wire                        cast_valid_i_2_23,
    output      wire                        cast_ready_o_2_23,

    output      wire        [`DW-1:0]       cast_data_o_2_23,
    output      wire                        cast_valid_o_2_23,
    input       wire                        cast_ready_i_2_23,

    input       wire        [`DW-1:0]       cast_data_i_2_24,
    input       wire                        cast_valid_i_2_24,
    output      wire                        cast_ready_o_2_24,

    output      wire        [`DW-1:0]       cast_data_o_2_24,
    output      wire                        cast_valid_o_2_24,
    input       wire                        cast_ready_i_2_24,

    input       wire        [`DW-1:0]       cast_data_i_3_0,
    input       wire                        cast_valid_i_3_0,
    output      wire                        cast_ready_o_3_0,

    output      wire        [`DW-1:0]       cast_data_o_3_0,
    output      wire                        cast_valid_o_3_0,
    input       wire                        cast_ready_i_3_0,

    input       wire        [`DW-1:0]       cast_data_i_3_1,
    input       wire                        cast_valid_i_3_1,
    output      wire                        cast_ready_o_3_1,

    output      wire        [`DW-1:0]       cast_data_o_3_1,
    output      wire                        cast_valid_o_3_1,
    input       wire                        cast_ready_i_3_1,

    input       wire        [`DW-1:0]       cast_data_i_3_2,
    input       wire                        cast_valid_i_3_2,
    output      wire                        cast_ready_o_3_2,

    output      wire        [`DW-1:0]       cast_data_o_3_2,
    output      wire                        cast_valid_o_3_2,
    input       wire                        cast_ready_i_3_2,

    input       wire        [`DW-1:0]       cast_data_i_3_3,
    input       wire                        cast_valid_i_3_3,
    output      wire                        cast_ready_o_3_3,

    output      wire        [`DW-1:0]       cast_data_o_3_3,
    output      wire                        cast_valid_o_3_3,
    input       wire                        cast_ready_i_3_3,

    input       wire        [`DW-1:0]       cast_data_i_3_4,
    input       wire                        cast_valid_i_3_4,
    output      wire                        cast_ready_o_3_4,

    output      wire        [`DW-1:0]       cast_data_o_3_4,
    output      wire                        cast_valid_o_3_4,
    input       wire                        cast_ready_i_3_4,

    input       wire        [`DW-1:0]       cast_data_i_3_5,
    input       wire                        cast_valid_i_3_5,
    output      wire                        cast_ready_o_3_5,

    output      wire        [`DW-1:0]       cast_data_o_3_5,
    output      wire                        cast_valid_o_3_5,
    input       wire                        cast_ready_i_3_5,

    input       wire        [`DW-1:0]       cast_data_i_3_6,
    input       wire                        cast_valid_i_3_6,
    output      wire                        cast_ready_o_3_6,

    output      wire        [`DW-1:0]       cast_data_o_3_6,
    output      wire                        cast_valid_o_3_6,
    input       wire                        cast_ready_i_3_6,

    input       wire        [`DW-1:0]       cast_data_i_3_7,
    input       wire                        cast_valid_i_3_7,
    output      wire                        cast_ready_o_3_7,

    output      wire        [`DW-1:0]       cast_data_o_3_7,
    output      wire                        cast_valid_o_3_7,
    input       wire                        cast_ready_i_3_7,

    input       wire        [`DW-1:0]       cast_data_i_3_8,
    input       wire                        cast_valid_i_3_8,
    output      wire                        cast_ready_o_3_8,

    output      wire        [`DW-1:0]       cast_data_o_3_8,
    output      wire                        cast_valid_o_3_8,
    input       wire                        cast_ready_i_3_8,

    input       wire        [`DW-1:0]       cast_data_i_3_9,
    input       wire                        cast_valid_i_3_9,
    output      wire                        cast_ready_o_3_9,

    output      wire        [`DW-1:0]       cast_data_o_3_9,
    output      wire                        cast_valid_o_3_9,
    input       wire                        cast_ready_i_3_9,

    input       wire        [`DW-1:0]       cast_data_i_3_10,
    input       wire                        cast_valid_i_3_10,
    output      wire                        cast_ready_o_3_10,

    output      wire        [`DW-1:0]       cast_data_o_3_10,
    output      wire                        cast_valid_o_3_10,
    input       wire                        cast_ready_i_3_10,

    input       wire        [`DW-1:0]       cast_data_i_3_11,
    input       wire                        cast_valid_i_3_11,
    output      wire                        cast_ready_o_3_11,

    output      wire        [`DW-1:0]       cast_data_o_3_11,
    output      wire                        cast_valid_o_3_11,
    input       wire                        cast_ready_i_3_11,

    input       wire        [`DW-1:0]       cast_data_i_3_12,
    input       wire                        cast_valid_i_3_12,
    output      wire                        cast_ready_o_3_12,

    output      wire        [`DW-1:0]       cast_data_o_3_12,
    output      wire                        cast_valid_o_3_12,
    input       wire                        cast_ready_i_3_12,

    input       wire        [`DW-1:0]       cast_data_i_3_13,
    input       wire                        cast_valid_i_3_13,
    output      wire                        cast_ready_o_3_13,

    output      wire        [`DW-1:0]       cast_data_o_3_13,
    output      wire                        cast_valid_o_3_13,
    input       wire                        cast_ready_i_3_13,

    input       wire        [`DW-1:0]       cast_data_i_3_14,
    input       wire                        cast_valid_i_3_14,
    output      wire                        cast_ready_o_3_14,

    output      wire        [`DW-1:0]       cast_data_o_3_14,
    output      wire                        cast_valid_o_3_14,
    input       wire                        cast_ready_i_3_14,

    input       wire        [`DW-1:0]       cast_data_i_3_15,
    input       wire                        cast_valid_i_3_15,
    output      wire                        cast_ready_o_3_15,

    output      wire        [`DW-1:0]       cast_data_o_3_15,
    output      wire                        cast_valid_o_3_15,
    input       wire                        cast_ready_i_3_15,

    input       wire        [`DW-1:0]       cast_data_i_3_16,
    input       wire                        cast_valid_i_3_16,
    output      wire                        cast_ready_o_3_16,

    output      wire        [`DW-1:0]       cast_data_o_3_16,
    output      wire                        cast_valid_o_3_16,
    input       wire                        cast_ready_i_3_16,

    input       wire        [`DW-1:0]       cast_data_i_3_17,
    input       wire                        cast_valid_i_3_17,
    output      wire                        cast_ready_o_3_17,

    output      wire        [`DW-1:0]       cast_data_o_3_17,
    output      wire                        cast_valid_o_3_17,
    input       wire                        cast_ready_i_3_17,

    input       wire        [`DW-1:0]       cast_data_i_3_18,
    input       wire                        cast_valid_i_3_18,
    output      wire                        cast_ready_o_3_18,

    output      wire        [`DW-1:0]       cast_data_o_3_18,
    output      wire                        cast_valid_o_3_18,
    input       wire                        cast_ready_i_3_18,

    input       wire        [`DW-1:0]       cast_data_i_3_19,
    input       wire                        cast_valid_i_3_19,
    output      wire                        cast_ready_o_3_19,

    output      wire        [`DW-1:0]       cast_data_o_3_19,
    output      wire                        cast_valid_o_3_19,
    input       wire                        cast_ready_i_3_19,

    input       wire        [`DW-1:0]       cast_data_i_3_20,
    input       wire                        cast_valid_i_3_20,
    output      wire                        cast_ready_o_3_20,

    output      wire        [`DW-1:0]       cast_data_o_3_20,
    output      wire                        cast_valid_o_3_20,
    input       wire                        cast_ready_i_3_20,

    input       wire        [`DW-1:0]       cast_data_i_3_21,
    input       wire                        cast_valid_i_3_21,
    output      wire                        cast_ready_o_3_21,

    output      wire        [`DW-1:0]       cast_data_o_3_21,
    output      wire                        cast_valid_o_3_21,
    input       wire                        cast_ready_i_3_21,

    input       wire        [`DW-1:0]       cast_data_i_3_22,
    input       wire                        cast_valid_i_3_22,
    output      wire                        cast_ready_o_3_22,

    output      wire        [`DW-1:0]       cast_data_o_3_22,
    output      wire                        cast_valid_o_3_22,
    input       wire                        cast_ready_i_3_22,

    input       wire        [`DW-1:0]       cast_data_i_3_23,
    input       wire                        cast_valid_i_3_23,
    output      wire                        cast_ready_o_3_23,

    output      wire        [`DW-1:0]       cast_data_o_3_23,
    output      wire                        cast_valid_o_3_23,
    input       wire                        cast_ready_i_3_23,

    input       wire        [`DW-1:0]       cast_data_i_3_24,
    input       wire                        cast_valid_i_3_24,
    output      wire                        cast_ready_o_3_24,

    output      wire        [`DW-1:0]       cast_data_o_3_24,
    output      wire                        cast_valid_o_3_24,
    input       wire                        cast_ready_i_3_24,

    input       wire        [`DW-1:0]       cast_data_i_4_0,
    input       wire                        cast_valid_i_4_0,
    output      wire                        cast_ready_o_4_0,

    output      wire        [`DW-1:0]       cast_data_o_4_0,
    output      wire                        cast_valid_o_4_0,
    input       wire                        cast_ready_i_4_0,

    input       wire        [`DW-1:0]       cast_data_i_4_1,
    input       wire                        cast_valid_i_4_1,
    output      wire                        cast_ready_o_4_1,

    output      wire        [`DW-1:0]       cast_data_o_4_1,
    output      wire                        cast_valid_o_4_1,
    input       wire                        cast_ready_i_4_1,

    input       wire        [`DW-1:0]       cast_data_i_4_2,
    input       wire                        cast_valid_i_4_2,
    output      wire                        cast_ready_o_4_2,

    output      wire        [`DW-1:0]       cast_data_o_4_2,
    output      wire                        cast_valid_o_4_2,
    input       wire                        cast_ready_i_4_2,

    input       wire        [`DW-1:0]       cast_data_i_4_3,
    input       wire                        cast_valid_i_4_3,
    output      wire                        cast_ready_o_4_3,

    output      wire        [`DW-1:0]       cast_data_o_4_3,
    output      wire                        cast_valid_o_4_3,
    input       wire                        cast_ready_i_4_3,

    input       wire        [`DW-1:0]       cast_data_i_4_4,
    input       wire                        cast_valid_i_4_4,
    output      wire                        cast_ready_o_4_4,

    output      wire        [`DW-1:0]       cast_data_o_4_4,
    output      wire                        cast_valid_o_4_4,
    input       wire                        cast_ready_i_4_4,

    input       wire        [`DW-1:0]       cast_data_i_4_5,
    input       wire                        cast_valid_i_4_5,
    output      wire                        cast_ready_o_4_5,

    output      wire        [`DW-1:0]       cast_data_o_4_5,
    output      wire                        cast_valid_o_4_5,
    input       wire                        cast_ready_i_4_5,

    input       wire        [`DW-1:0]       cast_data_i_4_6,
    input       wire                        cast_valid_i_4_6,
    output      wire                        cast_ready_o_4_6,

    output      wire        [`DW-1:0]       cast_data_o_4_6,
    output      wire                        cast_valid_o_4_6,
    input       wire                        cast_ready_i_4_6,

    input       wire        [`DW-1:0]       cast_data_i_4_7,
    input       wire                        cast_valid_i_4_7,
    output      wire                        cast_ready_o_4_7,

    output      wire        [`DW-1:0]       cast_data_o_4_7,
    output      wire                        cast_valid_o_4_7,
    input       wire                        cast_ready_i_4_7,

    input       wire        [`DW-1:0]       cast_data_i_4_8,
    input       wire                        cast_valid_i_4_8,
    output      wire                        cast_ready_o_4_8,

    output      wire        [`DW-1:0]       cast_data_o_4_8,
    output      wire                        cast_valid_o_4_8,
    input       wire                        cast_ready_i_4_8,

    input       wire        [`DW-1:0]       cast_data_i_4_9,
    input       wire                        cast_valid_i_4_9,
    output      wire                        cast_ready_o_4_9,

    output      wire        [`DW-1:0]       cast_data_o_4_9,
    output      wire                        cast_valid_o_4_9,
    input       wire                        cast_ready_i_4_9,

    input       wire        [`DW-1:0]       cast_data_i_4_10,
    input       wire                        cast_valid_i_4_10,
    output      wire                        cast_ready_o_4_10,

    output      wire        [`DW-1:0]       cast_data_o_4_10,
    output      wire                        cast_valid_o_4_10,
    input       wire                        cast_ready_i_4_10,

    input       wire        [`DW-1:0]       cast_data_i_4_11,
    input       wire                        cast_valid_i_4_11,
    output      wire                        cast_ready_o_4_11,

    output      wire        [`DW-1:0]       cast_data_o_4_11,
    output      wire                        cast_valid_o_4_11,
    input       wire                        cast_ready_i_4_11,

    input       wire        [`DW-1:0]       cast_data_i_4_12,
    input       wire                        cast_valid_i_4_12,
    output      wire                        cast_ready_o_4_12,

    output      wire        [`DW-1:0]       cast_data_o_4_12,
    output      wire                        cast_valid_o_4_12,
    input       wire                        cast_ready_i_4_12,

    input       wire        [`DW-1:0]       cast_data_i_4_13,
    input       wire                        cast_valid_i_4_13,
    output      wire                        cast_ready_o_4_13,

    output      wire        [`DW-1:0]       cast_data_o_4_13,
    output      wire                        cast_valid_o_4_13,
    input       wire                        cast_ready_i_4_13,

    input       wire        [`DW-1:0]       cast_data_i_4_14,
    input       wire                        cast_valid_i_4_14,
    output      wire                        cast_ready_o_4_14,

    output      wire        [`DW-1:0]       cast_data_o_4_14,
    output      wire                        cast_valid_o_4_14,
    input       wire                        cast_ready_i_4_14,

    input       wire        [`DW-1:0]       cast_data_i_4_15,
    input       wire                        cast_valid_i_4_15,
    output      wire                        cast_ready_o_4_15,

    output      wire        [`DW-1:0]       cast_data_o_4_15,
    output      wire                        cast_valid_o_4_15,
    input       wire                        cast_ready_i_4_15,

    input       wire        [`DW-1:0]       cast_data_i_4_16,
    input       wire                        cast_valid_i_4_16,
    output      wire                        cast_ready_o_4_16,

    output      wire        [`DW-1:0]       cast_data_o_4_16,
    output      wire                        cast_valid_o_4_16,
    input       wire                        cast_ready_i_4_16,

    input       wire        [`DW-1:0]       cast_data_i_4_17,
    input       wire                        cast_valid_i_4_17,
    output      wire                        cast_ready_o_4_17,

    output      wire        [`DW-1:0]       cast_data_o_4_17,
    output      wire                        cast_valid_o_4_17,
    input       wire                        cast_ready_i_4_17,

    input       wire        [`DW-1:0]       cast_data_i_4_18,
    input       wire                        cast_valid_i_4_18,
    output      wire                        cast_ready_o_4_18,

    output      wire        [`DW-1:0]       cast_data_o_4_18,
    output      wire                        cast_valid_o_4_18,
    input       wire                        cast_ready_i_4_18,

    input       wire        [`DW-1:0]       cast_data_i_4_19,
    input       wire                        cast_valid_i_4_19,
    output      wire                        cast_ready_o_4_19,

    output      wire        [`DW-1:0]       cast_data_o_4_19,
    output      wire                        cast_valid_o_4_19,
    input       wire                        cast_ready_i_4_19,

    input       wire        [`DW-1:0]       cast_data_i_4_20,
    input       wire                        cast_valid_i_4_20,
    output      wire                        cast_ready_o_4_20,

    output      wire        [`DW-1:0]       cast_data_o_4_20,
    output      wire                        cast_valid_o_4_20,
    input       wire                        cast_ready_i_4_20,

    input       wire        [`DW-1:0]       cast_data_i_4_21,
    input       wire                        cast_valid_i_4_21,
    output      wire                        cast_ready_o_4_21,

    output      wire        [`DW-1:0]       cast_data_o_4_21,
    output      wire                        cast_valid_o_4_21,
    input       wire                        cast_ready_i_4_21,

    input       wire        [`DW-1:0]       cast_data_i_4_22,
    input       wire                        cast_valid_i_4_22,
    output      wire                        cast_ready_o_4_22,

    output      wire        [`DW-1:0]       cast_data_o_4_22,
    output      wire                        cast_valid_o_4_22,
    input       wire                        cast_ready_i_4_22,

    input       wire        [`DW-1:0]       cast_data_i_4_23,
    input       wire                        cast_valid_i_4_23,
    output      wire                        cast_ready_o_4_23,

    output      wire        [`DW-1:0]       cast_data_o_4_23,
    output      wire                        cast_valid_o_4_23,
    input       wire                        cast_ready_i_4_23,

    input       wire        [`DW-1:0]       cast_data_i_4_24,
    input       wire                        cast_valid_i_4_24,
    output      wire                        cast_ready_o_4_24,

    output      wire        [`DW-1:0]       cast_data_o_4_24,
    output      wire                        cast_valid_o_4_24,
    input       wire                        cast_ready_i_4_24,

    input       wire        [`DW-1:0]       cast_data_i_5_0,
    input       wire                        cast_valid_i_5_0,
    output      wire                        cast_ready_o_5_0,

    output      wire        [`DW-1:0]       cast_data_o_5_0,
    output      wire                        cast_valid_o_5_0,
    input       wire                        cast_ready_i_5_0,

    input       wire        [`DW-1:0]       cast_data_i_5_1,
    input       wire                        cast_valid_i_5_1,
    output      wire                        cast_ready_o_5_1,

    output      wire        [`DW-1:0]       cast_data_o_5_1,
    output      wire                        cast_valid_o_5_1,
    input       wire                        cast_ready_i_5_1,

    input       wire        [`DW-1:0]       cast_data_i_5_2,
    input       wire                        cast_valid_i_5_2,
    output      wire                        cast_ready_o_5_2,

    output      wire        [`DW-1:0]       cast_data_o_5_2,
    output      wire                        cast_valid_o_5_2,
    input       wire                        cast_ready_i_5_2,

    input       wire        [`DW-1:0]       cast_data_i_5_3,
    input       wire                        cast_valid_i_5_3,
    output      wire                        cast_ready_o_5_3,

    output      wire        [`DW-1:0]       cast_data_o_5_3,
    output      wire                        cast_valid_o_5_3,
    input       wire                        cast_ready_i_5_3,

    input       wire        [`DW-1:0]       cast_data_i_5_4,
    input       wire                        cast_valid_i_5_4,
    output      wire                        cast_ready_o_5_4,

    output      wire        [`DW-1:0]       cast_data_o_5_4,
    output      wire                        cast_valid_o_5_4,
    input       wire                        cast_ready_i_5_4,

    input       wire        [`DW-1:0]       cast_data_i_5_5,
    input       wire                        cast_valid_i_5_5,
    output      wire                        cast_ready_o_5_5,

    output      wire        [`DW-1:0]       cast_data_o_5_5,
    output      wire                        cast_valid_o_5_5,
    input       wire                        cast_ready_i_5_5,

    input       wire        [`DW-1:0]       cast_data_i_5_6,
    input       wire                        cast_valid_i_5_6,
    output      wire                        cast_ready_o_5_6,

    output      wire        [`DW-1:0]       cast_data_o_5_6,
    output      wire                        cast_valid_o_5_6,
    input       wire                        cast_ready_i_5_6,

    input       wire        [`DW-1:0]       cast_data_i_5_7,
    input       wire                        cast_valid_i_5_7,
    output      wire                        cast_ready_o_5_7,

    output      wire        [`DW-1:0]       cast_data_o_5_7,
    output      wire                        cast_valid_o_5_7,
    input       wire                        cast_ready_i_5_7,

    input       wire        [`DW-1:0]       cast_data_i_5_8,
    input       wire                        cast_valid_i_5_8,
    output      wire                        cast_ready_o_5_8,

    output      wire        [`DW-1:0]       cast_data_o_5_8,
    output      wire                        cast_valid_o_5_8,
    input       wire                        cast_ready_i_5_8,

    input       wire        [`DW-1:0]       cast_data_i_5_9,
    input       wire                        cast_valid_i_5_9,
    output      wire                        cast_ready_o_5_9,

    output      wire        [`DW-1:0]       cast_data_o_5_9,
    output      wire                        cast_valid_o_5_9,
    input       wire                        cast_ready_i_5_9,

    input       wire        [`DW-1:0]       cast_data_i_5_10,
    input       wire                        cast_valid_i_5_10,
    output      wire                        cast_ready_o_5_10,

    output      wire        [`DW-1:0]       cast_data_o_5_10,
    output      wire                        cast_valid_o_5_10,
    input       wire                        cast_ready_i_5_10,

    input       wire        [`DW-1:0]       cast_data_i_5_11,
    input       wire                        cast_valid_i_5_11,
    output      wire                        cast_ready_o_5_11,

    output      wire        [`DW-1:0]       cast_data_o_5_11,
    output      wire                        cast_valid_o_5_11,
    input       wire                        cast_ready_i_5_11,

    input       wire        [`DW-1:0]       cast_data_i_5_12,
    input       wire                        cast_valid_i_5_12,
    output      wire                        cast_ready_o_5_12,

    output      wire        [`DW-1:0]       cast_data_o_5_12,
    output      wire                        cast_valid_o_5_12,
    input       wire                        cast_ready_i_5_12,

    input       wire        [`DW-1:0]       cast_data_i_5_13,
    input       wire                        cast_valid_i_5_13,
    output      wire                        cast_ready_o_5_13,

    output      wire        [`DW-1:0]       cast_data_o_5_13,
    output      wire                        cast_valid_o_5_13,
    input       wire                        cast_ready_i_5_13,

    input       wire        [`DW-1:0]       cast_data_i_5_14,
    input       wire                        cast_valid_i_5_14,
    output      wire                        cast_ready_o_5_14,

    output      wire        [`DW-1:0]       cast_data_o_5_14,
    output      wire                        cast_valid_o_5_14,
    input       wire                        cast_ready_i_5_14,

    input       wire        [`DW-1:0]       cast_data_i_5_15,
    input       wire                        cast_valid_i_5_15,
    output      wire                        cast_ready_o_5_15,

    output      wire        [`DW-1:0]       cast_data_o_5_15,
    output      wire                        cast_valid_o_5_15,
    input       wire                        cast_ready_i_5_15,

    input       wire        [`DW-1:0]       cast_data_i_5_16,
    input       wire                        cast_valid_i_5_16,
    output      wire                        cast_ready_o_5_16,

    output      wire        [`DW-1:0]       cast_data_o_5_16,
    output      wire                        cast_valid_o_5_16,
    input       wire                        cast_ready_i_5_16,

    input       wire        [`DW-1:0]       cast_data_i_5_17,
    input       wire                        cast_valid_i_5_17,
    output      wire                        cast_ready_o_5_17,

    output      wire        [`DW-1:0]       cast_data_o_5_17,
    output      wire                        cast_valid_o_5_17,
    input       wire                        cast_ready_i_5_17,

    input       wire        [`DW-1:0]       cast_data_i_5_18,
    input       wire                        cast_valid_i_5_18,
    output      wire                        cast_ready_o_5_18,

    output      wire        [`DW-1:0]       cast_data_o_5_18,
    output      wire                        cast_valid_o_5_18,
    input       wire                        cast_ready_i_5_18,

    input       wire        [`DW-1:0]       cast_data_i_5_19,
    input       wire                        cast_valid_i_5_19,
    output      wire                        cast_ready_o_5_19,

    output      wire        [`DW-1:0]       cast_data_o_5_19,
    output      wire                        cast_valid_o_5_19,
    input       wire                        cast_ready_i_5_19,

    input       wire        [`DW-1:0]       cast_data_i_5_20,
    input       wire                        cast_valid_i_5_20,
    output      wire                        cast_ready_o_5_20,

    output      wire        [`DW-1:0]       cast_data_o_5_20,
    output      wire                        cast_valid_o_5_20,
    input       wire                        cast_ready_i_5_20,

    input       wire        [`DW-1:0]       cast_data_i_5_21,
    input       wire                        cast_valid_i_5_21,
    output      wire                        cast_ready_o_5_21,

    output      wire        [`DW-1:0]       cast_data_o_5_21,
    output      wire                        cast_valid_o_5_21,
    input       wire                        cast_ready_i_5_21,

    input       wire        [`DW-1:0]       cast_data_i_5_22,
    input       wire                        cast_valid_i_5_22,
    output      wire                        cast_ready_o_5_22,

    output      wire        [`DW-1:0]       cast_data_o_5_22,
    output      wire                        cast_valid_o_5_22,
    input       wire                        cast_ready_i_5_22,

    input       wire        [`DW-1:0]       cast_data_i_5_23,
    input       wire                        cast_valid_i_5_23,
    output      wire                        cast_ready_o_5_23,

    output      wire        [`DW-1:0]       cast_data_o_5_23,
    output      wire                        cast_valid_o_5_23,
    input       wire                        cast_ready_i_5_23,

    input       wire        [`DW-1:0]       cast_data_i_5_24,
    input       wire                        cast_valid_i_5_24,
    output      wire                        cast_ready_o_5_24,

    output      wire        [`DW-1:0]       cast_data_o_5_24,
    output      wire                        cast_valid_o_5_24,
    input       wire                        cast_ready_i_5_24,

    input       wire        [`DW-1:0]       cast_data_i_6_0,
    input       wire                        cast_valid_i_6_0,
    output      wire                        cast_ready_o_6_0,

    output      wire        [`DW-1:0]       cast_data_o_6_0,
    output      wire                        cast_valid_o_6_0,
    input       wire                        cast_ready_i_6_0,

    input       wire        [`DW-1:0]       cast_data_i_6_1,
    input       wire                        cast_valid_i_6_1,
    output      wire                        cast_ready_o_6_1,

    output      wire        [`DW-1:0]       cast_data_o_6_1,
    output      wire                        cast_valid_o_6_1,
    input       wire                        cast_ready_i_6_1,

    input       wire        [`DW-1:0]       cast_data_i_6_2,
    input       wire                        cast_valid_i_6_2,
    output      wire                        cast_ready_o_6_2,

    output      wire        [`DW-1:0]       cast_data_o_6_2,
    output      wire                        cast_valid_o_6_2,
    input       wire                        cast_ready_i_6_2,

    input       wire        [`DW-1:0]       cast_data_i_6_3,
    input       wire                        cast_valid_i_6_3,
    output      wire                        cast_ready_o_6_3,

    output      wire        [`DW-1:0]       cast_data_o_6_3,
    output      wire                        cast_valid_o_6_3,
    input       wire                        cast_ready_i_6_3,

    input       wire        [`DW-1:0]       cast_data_i_6_4,
    input       wire                        cast_valid_i_6_4,
    output      wire                        cast_ready_o_6_4,

    output      wire        [`DW-1:0]       cast_data_o_6_4,
    output      wire                        cast_valid_o_6_4,
    input       wire                        cast_ready_i_6_4,

    input       wire        [`DW-1:0]       cast_data_i_6_5,
    input       wire                        cast_valid_i_6_5,
    output      wire                        cast_ready_o_6_5,

    output      wire        [`DW-1:0]       cast_data_o_6_5,
    output      wire                        cast_valid_o_6_5,
    input       wire                        cast_ready_i_6_5,

    input       wire        [`DW-1:0]       cast_data_i_6_6,
    input       wire                        cast_valid_i_6_6,
    output      wire                        cast_ready_o_6_6,

    output      wire        [`DW-1:0]       cast_data_o_6_6,
    output      wire                        cast_valid_o_6_6,
    input       wire                        cast_ready_i_6_6,

    input       wire        [`DW-1:0]       cast_data_i_6_7,
    input       wire                        cast_valid_i_6_7,
    output      wire                        cast_ready_o_6_7,

    output      wire        [`DW-1:0]       cast_data_o_6_7,
    output      wire                        cast_valid_o_6_7,
    input       wire                        cast_ready_i_6_7,

    input       wire        [`DW-1:0]       cast_data_i_6_8,
    input       wire                        cast_valid_i_6_8,
    output      wire                        cast_ready_o_6_8,

    output      wire        [`DW-1:0]       cast_data_o_6_8,
    output      wire                        cast_valid_o_6_8,
    input       wire                        cast_ready_i_6_8,

    input       wire        [`DW-1:0]       cast_data_i_6_9,
    input       wire                        cast_valid_i_6_9,
    output      wire                        cast_ready_o_6_9,

    output      wire        [`DW-1:0]       cast_data_o_6_9,
    output      wire                        cast_valid_o_6_9,
    input       wire                        cast_ready_i_6_9,

    input       wire        [`DW-1:0]       cast_data_i_6_10,
    input       wire                        cast_valid_i_6_10,
    output      wire                        cast_ready_o_6_10,

    output      wire        [`DW-1:0]       cast_data_o_6_10,
    output      wire                        cast_valid_o_6_10,
    input       wire                        cast_ready_i_6_10,

    input       wire        [`DW-1:0]       cast_data_i_6_11,
    input       wire                        cast_valid_i_6_11,
    output      wire                        cast_ready_o_6_11,

    output      wire        [`DW-1:0]       cast_data_o_6_11,
    output      wire                        cast_valid_o_6_11,
    input       wire                        cast_ready_i_6_11,

    input       wire        [`DW-1:0]       cast_data_i_6_12,
    input       wire                        cast_valid_i_6_12,
    output      wire                        cast_ready_o_6_12,

    output      wire        [`DW-1:0]       cast_data_o_6_12,
    output      wire                        cast_valid_o_6_12,
    input       wire                        cast_ready_i_6_12,

    input       wire        [`DW-1:0]       cast_data_i_6_13,
    input       wire                        cast_valid_i_6_13,
    output      wire                        cast_ready_o_6_13,

    output      wire        [`DW-1:0]       cast_data_o_6_13,
    output      wire                        cast_valid_o_6_13,
    input       wire                        cast_ready_i_6_13,

    input       wire        [`DW-1:0]       cast_data_i_6_14,
    input       wire                        cast_valid_i_6_14,
    output      wire                        cast_ready_o_6_14,

    output      wire        [`DW-1:0]       cast_data_o_6_14,
    output      wire                        cast_valid_o_6_14,
    input       wire                        cast_ready_i_6_14,

    input       wire        [`DW-1:0]       cast_data_i_6_15,
    input       wire                        cast_valid_i_6_15,
    output      wire                        cast_ready_o_6_15,

    output      wire        [`DW-1:0]       cast_data_o_6_15,
    output      wire                        cast_valid_o_6_15,
    input       wire                        cast_ready_i_6_15,

    input       wire        [`DW-1:0]       cast_data_i_6_16,
    input       wire                        cast_valid_i_6_16,
    output      wire                        cast_ready_o_6_16,

    output      wire        [`DW-1:0]       cast_data_o_6_16,
    output      wire                        cast_valid_o_6_16,
    input       wire                        cast_ready_i_6_16,

    input       wire        [`DW-1:0]       cast_data_i_6_17,
    input       wire                        cast_valid_i_6_17,
    output      wire                        cast_ready_o_6_17,

    output      wire        [`DW-1:0]       cast_data_o_6_17,
    output      wire                        cast_valid_o_6_17,
    input       wire                        cast_ready_i_6_17,

    input       wire        [`DW-1:0]       cast_data_i_6_18,
    input       wire                        cast_valid_i_6_18,
    output      wire                        cast_ready_o_6_18,

    output      wire        [`DW-1:0]       cast_data_o_6_18,
    output      wire                        cast_valid_o_6_18,
    input       wire                        cast_ready_i_6_18,

    input       wire        [`DW-1:0]       cast_data_i_6_19,
    input       wire                        cast_valid_i_6_19,
    output      wire                        cast_ready_o_6_19,

    output      wire        [`DW-1:0]       cast_data_o_6_19,
    output      wire                        cast_valid_o_6_19,
    input       wire                        cast_ready_i_6_19,

    input       wire        [`DW-1:0]       cast_data_i_6_20,
    input       wire                        cast_valid_i_6_20,
    output      wire                        cast_ready_o_6_20,

    output      wire        [`DW-1:0]       cast_data_o_6_20,
    output      wire                        cast_valid_o_6_20,
    input       wire                        cast_ready_i_6_20,

    input       wire        [`DW-1:0]       cast_data_i_6_21,
    input       wire                        cast_valid_i_6_21,
    output      wire                        cast_ready_o_6_21,

    output      wire        [`DW-1:0]       cast_data_o_6_21,
    output      wire                        cast_valid_o_6_21,
    input       wire                        cast_ready_i_6_21,

    input       wire        [`DW-1:0]       cast_data_i_6_22,
    input       wire                        cast_valid_i_6_22,
    output      wire                        cast_ready_o_6_22,

    output      wire        [`DW-1:0]       cast_data_o_6_22,
    output      wire                        cast_valid_o_6_22,
    input       wire                        cast_ready_i_6_22,

    input       wire        [`DW-1:0]       cast_data_i_6_23,
    input       wire                        cast_valid_i_6_23,
    output      wire                        cast_ready_o_6_23,

    output      wire        [`DW-1:0]       cast_data_o_6_23,
    output      wire                        cast_valid_o_6_23,
    input       wire                        cast_ready_i_6_23,

    input       wire        [`DW-1:0]       cast_data_i_6_24,
    input       wire                        cast_valid_i_6_24,
    output      wire                        cast_ready_o_6_24,

    output      wire        [`DW-1:0]       cast_data_o_6_24,
    output      wire                        cast_valid_o_6_24,
    input       wire                        cast_ready_i_6_24,

    input       wire        [`DW-1:0]       cast_data_i_7_0,
    input       wire                        cast_valid_i_7_0,
    output      wire                        cast_ready_o_7_0,

    output      wire        [`DW-1:0]       cast_data_o_7_0,
    output      wire                        cast_valid_o_7_0,
    input       wire                        cast_ready_i_7_0,

    input       wire        [`DW-1:0]       cast_data_i_7_1,
    input       wire                        cast_valid_i_7_1,
    output      wire                        cast_ready_o_7_1,

    output      wire        [`DW-1:0]       cast_data_o_7_1,
    output      wire                        cast_valid_o_7_1,
    input       wire                        cast_ready_i_7_1,

    input       wire        [`DW-1:0]       cast_data_i_7_2,
    input       wire                        cast_valid_i_7_2,
    output      wire                        cast_ready_o_7_2,

    output      wire        [`DW-1:0]       cast_data_o_7_2,
    output      wire                        cast_valid_o_7_2,
    input       wire                        cast_ready_i_7_2,

    input       wire        [`DW-1:0]       cast_data_i_7_3,
    input       wire                        cast_valid_i_7_3,
    output      wire                        cast_ready_o_7_3,

    output      wire        [`DW-1:0]       cast_data_o_7_3,
    output      wire                        cast_valid_o_7_3,
    input       wire                        cast_ready_i_7_3,

    input       wire        [`DW-1:0]       cast_data_i_7_4,
    input       wire                        cast_valid_i_7_4,
    output      wire                        cast_ready_o_7_4,

    output      wire        [`DW-1:0]       cast_data_o_7_4,
    output      wire                        cast_valid_o_7_4,
    input       wire                        cast_ready_i_7_4,

    input       wire        [`DW-1:0]       cast_data_i_7_5,
    input       wire                        cast_valid_i_7_5,
    output      wire                        cast_ready_o_7_5,

    output      wire        [`DW-1:0]       cast_data_o_7_5,
    output      wire                        cast_valid_o_7_5,
    input       wire                        cast_ready_i_7_5,

    input       wire        [`DW-1:0]       cast_data_i_7_6,
    input       wire                        cast_valid_i_7_6,
    output      wire                        cast_ready_o_7_6,

    output      wire        [`DW-1:0]       cast_data_o_7_6,
    output      wire                        cast_valid_o_7_6,
    input       wire                        cast_ready_i_7_6,

    input       wire        [`DW-1:0]       cast_data_i_7_7,
    input       wire                        cast_valid_i_7_7,
    output      wire                        cast_ready_o_7_7,

    output      wire        [`DW-1:0]       cast_data_o_7_7,
    output      wire                        cast_valid_o_7_7,
    input       wire                        cast_ready_i_7_7,

    input       wire        [`DW-1:0]       cast_data_i_7_8,
    input       wire                        cast_valid_i_7_8,
    output      wire                        cast_ready_o_7_8,

    output      wire        [`DW-1:0]       cast_data_o_7_8,
    output      wire                        cast_valid_o_7_8,
    input       wire                        cast_ready_i_7_8,

    input       wire        [`DW-1:0]       cast_data_i_7_9,
    input       wire                        cast_valid_i_7_9,
    output      wire                        cast_ready_o_7_9,

    output      wire        [`DW-1:0]       cast_data_o_7_9,
    output      wire                        cast_valid_o_7_9,
    input       wire                        cast_ready_i_7_9,

    input       wire        [`DW-1:0]       cast_data_i_7_10,
    input       wire                        cast_valid_i_7_10,
    output      wire                        cast_ready_o_7_10,

    output      wire        [`DW-1:0]       cast_data_o_7_10,
    output      wire                        cast_valid_o_7_10,
    input       wire                        cast_ready_i_7_10,

    input       wire        [`DW-1:0]       cast_data_i_7_11,
    input       wire                        cast_valid_i_7_11,
    output      wire                        cast_ready_o_7_11,

    output      wire        [`DW-1:0]       cast_data_o_7_11,
    output      wire                        cast_valid_o_7_11,
    input       wire                        cast_ready_i_7_11,

    input       wire        [`DW-1:0]       cast_data_i_7_12,
    input       wire                        cast_valid_i_7_12,
    output      wire                        cast_ready_o_7_12,

    output      wire        [`DW-1:0]       cast_data_o_7_12,
    output      wire                        cast_valid_o_7_12,
    input       wire                        cast_ready_i_7_12,

    input       wire        [`DW-1:0]       cast_data_i_7_13,
    input       wire                        cast_valid_i_7_13,
    output      wire                        cast_ready_o_7_13,

    output      wire        [`DW-1:0]       cast_data_o_7_13,
    output      wire                        cast_valid_o_7_13,
    input       wire                        cast_ready_i_7_13,

    input       wire        [`DW-1:0]       cast_data_i_7_14,
    input       wire                        cast_valid_i_7_14,
    output      wire                        cast_ready_o_7_14,

    output      wire        [`DW-1:0]       cast_data_o_7_14,
    output      wire                        cast_valid_o_7_14,
    input       wire                        cast_ready_i_7_14,

    input       wire        [`DW-1:0]       cast_data_i_7_15,
    input       wire                        cast_valid_i_7_15,
    output      wire                        cast_ready_o_7_15,

    output      wire        [`DW-1:0]       cast_data_o_7_15,
    output      wire                        cast_valid_o_7_15,
    input       wire                        cast_ready_i_7_15,

    input       wire        [`DW-1:0]       cast_data_i_7_16,
    input       wire                        cast_valid_i_7_16,
    output      wire                        cast_ready_o_7_16,

    output      wire        [`DW-1:0]       cast_data_o_7_16,
    output      wire                        cast_valid_o_7_16,
    input       wire                        cast_ready_i_7_16,

    input       wire        [`DW-1:0]       cast_data_i_7_17,
    input       wire                        cast_valid_i_7_17,
    output      wire                        cast_ready_o_7_17,

    output      wire        [`DW-1:0]       cast_data_o_7_17,
    output      wire                        cast_valid_o_7_17,
    input       wire                        cast_ready_i_7_17,

    input       wire        [`DW-1:0]       cast_data_i_7_18,
    input       wire                        cast_valid_i_7_18,
    output      wire                        cast_ready_o_7_18,

    output      wire        [`DW-1:0]       cast_data_o_7_18,
    output      wire                        cast_valid_o_7_18,
    input       wire                        cast_ready_i_7_18,

    input       wire        [`DW-1:0]       cast_data_i_7_19,
    input       wire                        cast_valid_i_7_19,
    output      wire                        cast_ready_o_7_19,

    output      wire        [`DW-1:0]       cast_data_o_7_19,
    output      wire                        cast_valid_o_7_19,
    input       wire                        cast_ready_i_7_19,

    input       wire        [`DW-1:0]       cast_data_i_7_20,
    input       wire                        cast_valid_i_7_20,
    output      wire                        cast_ready_o_7_20,

    output      wire        [`DW-1:0]       cast_data_o_7_20,
    output      wire                        cast_valid_o_7_20,
    input       wire                        cast_ready_i_7_20,

    input       wire        [`DW-1:0]       cast_data_i_7_21,
    input       wire                        cast_valid_i_7_21,
    output      wire                        cast_ready_o_7_21,

    output      wire        [`DW-1:0]       cast_data_o_7_21,
    output      wire                        cast_valid_o_7_21,
    input       wire                        cast_ready_i_7_21,

    input       wire        [`DW-1:0]       cast_data_i_7_22,
    input       wire                        cast_valid_i_7_22,
    output      wire                        cast_ready_o_7_22,

    output      wire        [`DW-1:0]       cast_data_o_7_22,
    output      wire                        cast_valid_o_7_22,
    input       wire                        cast_ready_i_7_22,

    input       wire        [`DW-1:0]       cast_data_i_7_23,
    input       wire                        cast_valid_i_7_23,
    output      wire                        cast_ready_o_7_23,

    output      wire        [`DW-1:0]       cast_data_o_7_23,
    output      wire                        cast_valid_o_7_23,
    input       wire                        cast_ready_i_7_23,

    input       wire        [`DW-1:0]       cast_data_i_7_24,
    input       wire                        cast_valid_i_7_24,
    output      wire                        cast_ready_o_7_24,

    output      wire        [`DW-1:0]       cast_data_o_7_24,
    output      wire                        cast_valid_o_7_24,
    input       wire                        cast_ready_i_7_24,

    input       wire        [`DW-1:0]       cast_data_i_8_0,
    input       wire                        cast_valid_i_8_0,
    output      wire                        cast_ready_o_8_0,

    output      wire        [`DW-1:0]       cast_data_o_8_0,
    output      wire                        cast_valid_o_8_0,
    input       wire                        cast_ready_i_8_0,

    input       wire        [`DW-1:0]       cast_data_i_8_1,
    input       wire                        cast_valid_i_8_1,
    output      wire                        cast_ready_o_8_1,

    output      wire        [`DW-1:0]       cast_data_o_8_1,
    output      wire                        cast_valid_o_8_1,
    input       wire                        cast_ready_i_8_1,

    input       wire        [`DW-1:0]       cast_data_i_8_2,
    input       wire                        cast_valid_i_8_2,
    output      wire                        cast_ready_o_8_2,

    output      wire        [`DW-1:0]       cast_data_o_8_2,
    output      wire                        cast_valid_o_8_2,
    input       wire                        cast_ready_i_8_2,

    input       wire        [`DW-1:0]       cast_data_i_8_3,
    input       wire                        cast_valid_i_8_3,
    output      wire                        cast_ready_o_8_3,

    output      wire        [`DW-1:0]       cast_data_o_8_3,
    output      wire                        cast_valid_o_8_3,
    input       wire                        cast_ready_i_8_3,

    input       wire        [`DW-1:0]       cast_data_i_8_4,
    input       wire                        cast_valid_i_8_4,
    output      wire                        cast_ready_o_8_4,

    output      wire        [`DW-1:0]       cast_data_o_8_4,
    output      wire                        cast_valid_o_8_4,
    input       wire                        cast_ready_i_8_4,

    input       wire        [`DW-1:0]       cast_data_i_8_5,
    input       wire                        cast_valid_i_8_5,
    output      wire                        cast_ready_o_8_5,

    output      wire        [`DW-1:0]       cast_data_o_8_5,
    output      wire                        cast_valid_o_8_5,
    input       wire                        cast_ready_i_8_5,

    input       wire        [`DW-1:0]       cast_data_i_8_6,
    input       wire                        cast_valid_i_8_6,
    output      wire                        cast_ready_o_8_6,

    output      wire        [`DW-1:0]       cast_data_o_8_6,
    output      wire                        cast_valid_o_8_6,
    input       wire                        cast_ready_i_8_6,

    input       wire        [`DW-1:0]       cast_data_i_8_7,
    input       wire                        cast_valid_i_8_7,
    output      wire                        cast_ready_o_8_7,

    output      wire        [`DW-1:0]       cast_data_o_8_7,
    output      wire                        cast_valid_o_8_7,
    input       wire                        cast_ready_i_8_7,

    input       wire        [`DW-1:0]       cast_data_i_8_8,
    input       wire                        cast_valid_i_8_8,
    output      wire                        cast_ready_o_8_8,

    output      wire        [`DW-1:0]       cast_data_o_8_8,
    output      wire                        cast_valid_o_8_8,
    input       wire                        cast_ready_i_8_8,

    input       wire        [`DW-1:0]       cast_data_i_8_9,
    input       wire                        cast_valid_i_8_9,
    output      wire                        cast_ready_o_8_9,

    output      wire        [`DW-1:0]       cast_data_o_8_9,
    output      wire                        cast_valid_o_8_9,
    input       wire                        cast_ready_i_8_9,

    input       wire        [`DW-1:0]       cast_data_i_8_10,
    input       wire                        cast_valid_i_8_10,
    output      wire                        cast_ready_o_8_10,

    output      wire        [`DW-1:0]       cast_data_o_8_10,
    output      wire                        cast_valid_o_8_10,
    input       wire                        cast_ready_i_8_10,

    input       wire        [`DW-1:0]       cast_data_i_8_11,
    input       wire                        cast_valid_i_8_11,
    output      wire                        cast_ready_o_8_11,

    output      wire        [`DW-1:0]       cast_data_o_8_11,
    output      wire                        cast_valid_o_8_11,
    input       wire                        cast_ready_i_8_11,

    input       wire        [`DW-1:0]       cast_data_i_8_12,
    input       wire                        cast_valid_i_8_12,
    output      wire                        cast_ready_o_8_12,

    output      wire        [`DW-1:0]       cast_data_o_8_12,
    output      wire                        cast_valid_o_8_12,
    input       wire                        cast_ready_i_8_12,

    input       wire        [`DW-1:0]       cast_data_i_8_13,
    input       wire                        cast_valid_i_8_13,
    output      wire                        cast_ready_o_8_13,

    output      wire        [`DW-1:0]       cast_data_o_8_13,
    output      wire                        cast_valid_o_8_13,
    input       wire                        cast_ready_i_8_13,

    input       wire        [`DW-1:0]       cast_data_i_8_14,
    input       wire                        cast_valid_i_8_14,
    output      wire                        cast_ready_o_8_14,

    output      wire        [`DW-1:0]       cast_data_o_8_14,
    output      wire                        cast_valid_o_8_14,
    input       wire                        cast_ready_i_8_14,

    input       wire        [`DW-1:0]       cast_data_i_8_15,
    input       wire                        cast_valid_i_8_15,
    output      wire                        cast_ready_o_8_15,

    output      wire        [`DW-1:0]       cast_data_o_8_15,
    output      wire                        cast_valid_o_8_15,
    input       wire                        cast_ready_i_8_15,

    input       wire        [`DW-1:0]       cast_data_i_8_16,
    input       wire                        cast_valid_i_8_16,
    output      wire                        cast_ready_o_8_16,

    output      wire        [`DW-1:0]       cast_data_o_8_16,
    output      wire                        cast_valid_o_8_16,
    input       wire                        cast_ready_i_8_16,

    input       wire        [`DW-1:0]       cast_data_i_8_17,
    input       wire                        cast_valid_i_8_17,
    output      wire                        cast_ready_o_8_17,

    output      wire        [`DW-1:0]       cast_data_o_8_17,
    output      wire                        cast_valid_o_8_17,
    input       wire                        cast_ready_i_8_17,

    input       wire        [`DW-1:0]       cast_data_i_8_18,
    input       wire                        cast_valid_i_8_18,
    output      wire                        cast_ready_o_8_18,

    output      wire        [`DW-1:0]       cast_data_o_8_18,
    output      wire                        cast_valid_o_8_18,
    input       wire                        cast_ready_i_8_18,

    input       wire        [`DW-1:0]       cast_data_i_8_19,
    input       wire                        cast_valid_i_8_19,
    output      wire                        cast_ready_o_8_19,

    output      wire        [`DW-1:0]       cast_data_o_8_19,
    output      wire                        cast_valid_o_8_19,
    input       wire                        cast_ready_i_8_19,

    input       wire        [`DW-1:0]       cast_data_i_8_20,
    input       wire                        cast_valid_i_8_20,
    output      wire                        cast_ready_o_8_20,

    output      wire        [`DW-1:0]       cast_data_o_8_20,
    output      wire                        cast_valid_o_8_20,
    input       wire                        cast_ready_i_8_20,

    input       wire        [`DW-1:0]       cast_data_i_8_21,
    input       wire                        cast_valid_i_8_21,
    output      wire                        cast_ready_o_8_21,

    output      wire        [`DW-1:0]       cast_data_o_8_21,
    output      wire                        cast_valid_o_8_21,
    input       wire                        cast_ready_i_8_21,

    input       wire        [`DW-1:0]       cast_data_i_8_22,
    input       wire                        cast_valid_i_8_22,
    output      wire                        cast_ready_o_8_22,

    output      wire        [`DW-1:0]       cast_data_o_8_22,
    output      wire                        cast_valid_o_8_22,
    input       wire                        cast_ready_i_8_22,

    input       wire        [`DW-1:0]       cast_data_i_8_23,
    input       wire                        cast_valid_i_8_23,
    output      wire                        cast_ready_o_8_23,

    output      wire        [`DW-1:0]       cast_data_o_8_23,
    output      wire                        cast_valid_o_8_23,
    input       wire                        cast_ready_i_8_23,

    input       wire        [`DW-1:0]       cast_data_i_8_24,
    input       wire                        cast_valid_i_8_24,
    output      wire                        cast_ready_o_8_24,

    output      wire        [`DW-1:0]       cast_data_o_8_24,
    output      wire                        cast_valid_o_8_24,
    input       wire                        cast_ready_i_8_24,

    input       wire        [`DW-1:0]       cast_data_i_9_0,
    input       wire                        cast_valid_i_9_0,
    output      wire                        cast_ready_o_9_0,

    output      wire        [`DW-1:0]       cast_data_o_9_0,
    output      wire                        cast_valid_o_9_0,
    input       wire                        cast_ready_i_9_0,

    input       wire        [`DW-1:0]       cast_data_i_9_1,
    input       wire                        cast_valid_i_9_1,
    output      wire                        cast_ready_o_9_1,

    output      wire        [`DW-1:0]       cast_data_o_9_1,
    output      wire                        cast_valid_o_9_1,
    input       wire                        cast_ready_i_9_1,

    input       wire        [`DW-1:0]       cast_data_i_9_2,
    input       wire                        cast_valid_i_9_2,
    output      wire                        cast_ready_o_9_2,

    output      wire        [`DW-1:0]       cast_data_o_9_2,
    output      wire                        cast_valid_o_9_2,
    input       wire                        cast_ready_i_9_2,

    input       wire        [`DW-1:0]       cast_data_i_9_3,
    input       wire                        cast_valid_i_9_3,
    output      wire                        cast_ready_o_9_3,

    output      wire        [`DW-1:0]       cast_data_o_9_3,
    output      wire                        cast_valid_o_9_3,
    input       wire                        cast_ready_i_9_3,

    input       wire        [`DW-1:0]       cast_data_i_9_4,
    input       wire                        cast_valid_i_9_4,
    output      wire                        cast_ready_o_9_4,

    output      wire        [`DW-1:0]       cast_data_o_9_4,
    output      wire                        cast_valid_o_9_4,
    input       wire                        cast_ready_i_9_4,

    input       wire        [`DW-1:0]       cast_data_i_9_5,
    input       wire                        cast_valid_i_9_5,
    output      wire                        cast_ready_o_9_5,

    output      wire        [`DW-1:0]       cast_data_o_9_5,
    output      wire                        cast_valid_o_9_5,
    input       wire                        cast_ready_i_9_5,

    input       wire        [`DW-1:0]       cast_data_i_9_6,
    input       wire                        cast_valid_i_9_6,
    output      wire                        cast_ready_o_9_6,

    output      wire        [`DW-1:0]       cast_data_o_9_6,
    output      wire                        cast_valid_o_9_6,
    input       wire                        cast_ready_i_9_6,

    input       wire        [`DW-1:0]       cast_data_i_9_7,
    input       wire                        cast_valid_i_9_7,
    output      wire                        cast_ready_o_9_7,

    output      wire        [`DW-1:0]       cast_data_o_9_7,
    output      wire                        cast_valid_o_9_7,
    input       wire                        cast_ready_i_9_7,

    input       wire        [`DW-1:0]       cast_data_i_9_8,
    input       wire                        cast_valid_i_9_8,
    output      wire                        cast_ready_o_9_8,

    output      wire        [`DW-1:0]       cast_data_o_9_8,
    output      wire                        cast_valid_o_9_8,
    input       wire                        cast_ready_i_9_8,

    input       wire        [`DW-1:0]       cast_data_i_9_9,
    input       wire                        cast_valid_i_9_9,
    output      wire                        cast_ready_o_9_9,

    output      wire        [`DW-1:0]       cast_data_o_9_9,
    output      wire                        cast_valid_o_9_9,
    input       wire                        cast_ready_i_9_9,

    input       wire        [`DW-1:0]       cast_data_i_9_10,
    input       wire                        cast_valid_i_9_10,
    output      wire                        cast_ready_o_9_10,

    output      wire        [`DW-1:0]       cast_data_o_9_10,
    output      wire                        cast_valid_o_9_10,
    input       wire                        cast_ready_i_9_10,

    input       wire        [`DW-1:0]       cast_data_i_9_11,
    input       wire                        cast_valid_i_9_11,
    output      wire                        cast_ready_o_9_11,

    output      wire        [`DW-1:0]       cast_data_o_9_11,
    output      wire                        cast_valid_o_9_11,
    input       wire                        cast_ready_i_9_11,

    input       wire        [`DW-1:0]       cast_data_i_9_12,
    input       wire                        cast_valid_i_9_12,
    output      wire                        cast_ready_o_9_12,

    output      wire        [`DW-1:0]       cast_data_o_9_12,
    output      wire                        cast_valid_o_9_12,
    input       wire                        cast_ready_i_9_12,

    input       wire        [`DW-1:0]       cast_data_i_9_13,
    input       wire                        cast_valid_i_9_13,
    output      wire                        cast_ready_o_9_13,

    output      wire        [`DW-1:0]       cast_data_o_9_13,
    output      wire                        cast_valid_o_9_13,
    input       wire                        cast_ready_i_9_13,

    input       wire        [`DW-1:0]       cast_data_i_9_14,
    input       wire                        cast_valid_i_9_14,
    output      wire                        cast_ready_o_9_14,

    output      wire        [`DW-1:0]       cast_data_o_9_14,
    output      wire                        cast_valid_o_9_14,
    input       wire                        cast_ready_i_9_14,

    input       wire        [`DW-1:0]       cast_data_i_9_15,
    input       wire                        cast_valid_i_9_15,
    output      wire                        cast_ready_o_9_15,

    output      wire        [`DW-1:0]       cast_data_o_9_15,
    output      wire                        cast_valid_o_9_15,
    input       wire                        cast_ready_i_9_15,

    input       wire        [`DW-1:0]       cast_data_i_9_16,
    input       wire                        cast_valid_i_9_16,
    output      wire                        cast_ready_o_9_16,

    output      wire        [`DW-1:0]       cast_data_o_9_16,
    output      wire                        cast_valid_o_9_16,
    input       wire                        cast_ready_i_9_16,

    input       wire        [`DW-1:0]       cast_data_i_9_17,
    input       wire                        cast_valid_i_9_17,
    output      wire                        cast_ready_o_9_17,

    output      wire        [`DW-1:0]       cast_data_o_9_17,
    output      wire                        cast_valid_o_9_17,
    input       wire                        cast_ready_i_9_17,

    input       wire        [`DW-1:0]       cast_data_i_9_18,
    input       wire                        cast_valid_i_9_18,
    output      wire                        cast_ready_o_9_18,

    output      wire        [`DW-1:0]       cast_data_o_9_18,
    output      wire                        cast_valid_o_9_18,
    input       wire                        cast_ready_i_9_18,

    input       wire        [`DW-1:0]       cast_data_i_9_19,
    input       wire                        cast_valid_i_9_19,
    output      wire                        cast_ready_o_9_19,

    output      wire        [`DW-1:0]       cast_data_o_9_19,
    output      wire                        cast_valid_o_9_19,
    input       wire                        cast_ready_i_9_19,

    input       wire        [`DW-1:0]       cast_data_i_9_20,
    input       wire                        cast_valid_i_9_20,
    output      wire                        cast_ready_o_9_20,

    output      wire        [`DW-1:0]       cast_data_o_9_20,
    output      wire                        cast_valid_o_9_20,
    input       wire                        cast_ready_i_9_20,

    input       wire        [`DW-1:0]       cast_data_i_9_21,
    input       wire                        cast_valid_i_9_21,
    output      wire                        cast_ready_o_9_21,

    output      wire        [`DW-1:0]       cast_data_o_9_21,
    output      wire                        cast_valid_o_9_21,
    input       wire                        cast_ready_i_9_21,

    input       wire        [`DW-1:0]       cast_data_i_9_22,
    input       wire                        cast_valid_i_9_22,
    output      wire                        cast_ready_o_9_22,

    output      wire        [`DW-1:0]       cast_data_o_9_22,
    output      wire                        cast_valid_o_9_22,
    input       wire                        cast_ready_i_9_22,

    input       wire        [`DW-1:0]       cast_data_i_9_23,
    input       wire                        cast_valid_i_9_23,
    output      wire                        cast_ready_o_9_23,

    output      wire        [`DW-1:0]       cast_data_o_9_23,
    output      wire                        cast_valid_o_9_23,
    input       wire                        cast_ready_i_9_23,

    input       wire        [`DW-1:0]       cast_data_i_9_24,
    input       wire                        cast_valid_i_9_24,
    output      wire                        cast_ready_o_9_24,

    output      wire        [`DW-1:0]       cast_data_o_9_24,
    output      wire                        cast_valid_o_9_24,
    input       wire                        cast_ready_i_9_24,

    input       wire        [`DW-1:0]       merge_data_i_0_0,
    input       wire                        merge_valid_i_0_0,
    output      wire                        merge_ready_o_0_0,

    output      wire        [`DW-1:0]       merge_data_o_0_0,
    output      wire                        merge_valid_o_0_0,
    input       wire                        merge_ready_i_0_0,
    input       wire        [`DW-1:0]       merge_data_i_0_1,
    input       wire                        merge_valid_i_0_1,
    output      wire                        merge_ready_o_0_1,

    output      wire        [`DW-1:0]       merge_data_o_0_1,
    output      wire                        merge_valid_o_0_1,
    input       wire                        merge_ready_i_0_1,
    input       wire        [`DW-1:0]       merge_data_i_0_2,
    input       wire                        merge_valid_i_0_2,
    output      wire                        merge_ready_o_0_2,

    output      wire        [`DW-1:0]       merge_data_o_0_2,
    output      wire                        merge_valid_o_0_2,
    input       wire                        merge_ready_i_0_2,
    input       wire        [`DW-1:0]       merge_data_i_0_3,
    input       wire                        merge_valid_i_0_3,
    output      wire                        merge_ready_o_0_3,

    output      wire        [`DW-1:0]       merge_data_o_0_3,
    output      wire                        merge_valid_o_0_3,
    input       wire                        merge_ready_i_0_3,
    input       wire        [`DW-1:0]       merge_data_i_0_4,
    input       wire                        merge_valid_i_0_4,
    output      wire                        merge_ready_o_0_4,

    output      wire        [`DW-1:0]       merge_data_o_0_4,
    output      wire                        merge_valid_o_0_4,
    input       wire                        merge_ready_i_0_4,
    input       wire        [`DW-1:0]       merge_data_i_0_5,
    input       wire                        merge_valid_i_0_5,
    output      wire                        merge_ready_o_0_5,

    output      wire        [`DW-1:0]       merge_data_o_0_5,
    output      wire                        merge_valid_o_0_5,
    input       wire                        merge_ready_i_0_5,
    input       wire        [`DW-1:0]       merge_data_i_0_6,
    input       wire                        merge_valid_i_0_6,
    output      wire                        merge_ready_o_0_6,

    output      wire        [`DW-1:0]       merge_data_o_0_6,
    output      wire                        merge_valid_o_0_6,
    input       wire                        merge_ready_i_0_6,
    input       wire        [`DW-1:0]       merge_data_i_0_7,
    input       wire                        merge_valid_i_0_7,
    output      wire                        merge_ready_o_0_7,

    output      wire        [`DW-1:0]       merge_data_o_0_7,
    output      wire                        merge_valid_o_0_7,
    input       wire                        merge_ready_i_0_7,
    input       wire        [`DW-1:0]       merge_data_i_0_8,
    input       wire                        merge_valid_i_0_8,
    output      wire                        merge_ready_o_0_8,

    output      wire        [`DW-1:0]       merge_data_o_0_8,
    output      wire                        merge_valid_o_0_8,
    input       wire                        merge_ready_i_0_8,
    input       wire        [`DW-1:0]       merge_data_i_0_9,
    input       wire                        merge_valid_i_0_9,
    output      wire                        merge_ready_o_0_9,

    output      wire        [`DW-1:0]       merge_data_o_0_9,
    output      wire                        merge_valid_o_0_9,
    input       wire                        merge_ready_i_0_9,
    input       wire        [`DW-1:0]       merge_data_i_0_10,
    input       wire                        merge_valid_i_0_10,
    output      wire                        merge_ready_o_0_10,

    output      wire        [`DW-1:0]       merge_data_o_0_10,
    output      wire                        merge_valid_o_0_10,
    input       wire                        merge_ready_i_0_10,
    input       wire        [`DW-1:0]       merge_data_i_0_11,
    input       wire                        merge_valid_i_0_11,
    output      wire                        merge_ready_o_0_11,

    output      wire        [`DW-1:0]       merge_data_o_0_11,
    output      wire                        merge_valid_o_0_11,
    input       wire                        merge_ready_i_0_11,
    input       wire        [`DW-1:0]       merge_data_i_0_12,
    input       wire                        merge_valid_i_0_12,
    output      wire                        merge_ready_o_0_12,

    output      wire        [`DW-1:0]       merge_data_o_0_12,
    output      wire                        merge_valid_o_0_12,
    input       wire                        merge_ready_i_0_12,
    input       wire        [`DW-1:0]       merge_data_i_0_13,
    input       wire                        merge_valid_i_0_13,
    output      wire                        merge_ready_o_0_13,

    output      wire        [`DW-1:0]       merge_data_o_0_13,
    output      wire                        merge_valid_o_0_13,
    input       wire                        merge_ready_i_0_13,
    input       wire        [`DW-1:0]       merge_data_i_0_14,
    input       wire                        merge_valid_i_0_14,
    output      wire                        merge_ready_o_0_14,

    output      wire        [`DW-1:0]       merge_data_o_0_14,
    output      wire                        merge_valid_o_0_14,
    input       wire                        merge_ready_i_0_14,
    input       wire        [`DW-1:0]       merge_data_i_0_15,
    input       wire                        merge_valid_i_0_15,
    output      wire                        merge_ready_o_0_15,

    output      wire        [`DW-1:0]       merge_data_o_0_15,
    output      wire                        merge_valid_o_0_15,
    input       wire                        merge_ready_i_0_15,
    input       wire        [`DW-1:0]       merge_data_i_0_16,
    input       wire                        merge_valid_i_0_16,
    output      wire                        merge_ready_o_0_16,

    output      wire        [`DW-1:0]       merge_data_o_0_16,
    output      wire                        merge_valid_o_0_16,
    input       wire                        merge_ready_i_0_16,
    input       wire        [`DW-1:0]       merge_data_i_0_17,
    input       wire                        merge_valid_i_0_17,
    output      wire                        merge_ready_o_0_17,

    output      wire        [`DW-1:0]       merge_data_o_0_17,
    output      wire                        merge_valid_o_0_17,
    input       wire                        merge_ready_i_0_17,
    input       wire        [`DW-1:0]       merge_data_i_0_18,
    input       wire                        merge_valid_i_0_18,
    output      wire                        merge_ready_o_0_18,

    output      wire        [`DW-1:0]       merge_data_o_0_18,
    output      wire                        merge_valid_o_0_18,
    input       wire                        merge_ready_i_0_18,
    input       wire        [`DW-1:0]       merge_data_i_0_19,
    input       wire                        merge_valid_i_0_19,
    output      wire                        merge_ready_o_0_19,

    output      wire        [`DW-1:0]       merge_data_o_0_19,
    output      wire                        merge_valid_o_0_19,
    input       wire                        merge_ready_i_0_19,
    input       wire        [`DW-1:0]       merge_data_i_0_20,
    input       wire                        merge_valid_i_0_20,
    output      wire                        merge_ready_o_0_20,

    output      wire        [`DW-1:0]       merge_data_o_0_20,
    output      wire                        merge_valid_o_0_20,
    input       wire                        merge_ready_i_0_20,
    input       wire        [`DW-1:0]       merge_data_i_0_21,
    input       wire                        merge_valid_i_0_21,
    output      wire                        merge_ready_o_0_21,

    output      wire        [`DW-1:0]       merge_data_o_0_21,
    output      wire                        merge_valid_o_0_21,
    input       wire                        merge_ready_i_0_21,
    input       wire        [`DW-1:0]       merge_data_i_0_22,
    input       wire                        merge_valid_i_0_22,
    output      wire                        merge_ready_o_0_22,

    output      wire        [`DW-1:0]       merge_data_o_0_22,
    output      wire                        merge_valid_o_0_22,
    input       wire                        merge_ready_i_0_22,
    input       wire        [`DW-1:0]       merge_data_i_0_23,
    input       wire                        merge_valid_i_0_23,
    output      wire                        merge_ready_o_0_23,

    output      wire        [`DW-1:0]       merge_data_o_0_23,
    output      wire                        merge_valid_o_0_23,
    input       wire                        merge_ready_i_0_23,
    input       wire        [`DW-1:0]       merge_data_i_0_24,
    input       wire                        merge_valid_i_0_24,
    output      wire                        merge_ready_o_0_24,

    output      wire        [`DW-1:0]       merge_data_o_0_24,
    output      wire                        merge_valid_o_0_24,
    input       wire                        merge_ready_i_0_24,
    input       wire        [`DW-1:0]       merge_data_i_1_0,
    input       wire                        merge_valid_i_1_0,
    output      wire                        merge_ready_o_1_0,

    output      wire        [`DW-1:0]       merge_data_o_1_0,
    output      wire                        merge_valid_o_1_0,
    input       wire                        merge_ready_i_1_0,
    input       wire        [`DW-1:0]       merge_data_i_1_1,
    input       wire                        merge_valid_i_1_1,
    output      wire                        merge_ready_o_1_1,

    output      wire        [`DW-1:0]       merge_data_o_1_1,
    output      wire                        merge_valid_o_1_1,
    input       wire                        merge_ready_i_1_1,
    input       wire        [`DW-1:0]       merge_data_i_1_2,
    input       wire                        merge_valid_i_1_2,
    output      wire                        merge_ready_o_1_2,

    output      wire        [`DW-1:0]       merge_data_o_1_2,
    output      wire                        merge_valid_o_1_2,
    input       wire                        merge_ready_i_1_2,
    input       wire        [`DW-1:0]       merge_data_i_1_3,
    input       wire                        merge_valid_i_1_3,
    output      wire                        merge_ready_o_1_3,

    output      wire        [`DW-1:0]       merge_data_o_1_3,
    output      wire                        merge_valid_o_1_3,
    input       wire                        merge_ready_i_1_3,
    input       wire        [`DW-1:0]       merge_data_i_1_4,
    input       wire                        merge_valid_i_1_4,
    output      wire                        merge_ready_o_1_4,

    output      wire        [`DW-1:0]       merge_data_o_1_4,
    output      wire                        merge_valid_o_1_4,
    input       wire                        merge_ready_i_1_4,
    input       wire        [`DW-1:0]       merge_data_i_1_5,
    input       wire                        merge_valid_i_1_5,
    output      wire                        merge_ready_o_1_5,

    output      wire        [`DW-1:0]       merge_data_o_1_5,
    output      wire                        merge_valid_o_1_5,
    input       wire                        merge_ready_i_1_5,
    input       wire        [`DW-1:0]       merge_data_i_1_6,
    input       wire                        merge_valid_i_1_6,
    output      wire                        merge_ready_o_1_6,

    output      wire        [`DW-1:0]       merge_data_o_1_6,
    output      wire                        merge_valid_o_1_6,
    input       wire                        merge_ready_i_1_6,
    input       wire        [`DW-1:0]       merge_data_i_1_7,
    input       wire                        merge_valid_i_1_7,
    output      wire                        merge_ready_o_1_7,

    output      wire        [`DW-1:0]       merge_data_o_1_7,
    output      wire                        merge_valid_o_1_7,
    input       wire                        merge_ready_i_1_7,
    input       wire        [`DW-1:0]       merge_data_i_1_8,
    input       wire                        merge_valid_i_1_8,
    output      wire                        merge_ready_o_1_8,

    output      wire        [`DW-1:0]       merge_data_o_1_8,
    output      wire                        merge_valid_o_1_8,
    input       wire                        merge_ready_i_1_8,
    input       wire        [`DW-1:0]       merge_data_i_1_9,
    input       wire                        merge_valid_i_1_9,
    output      wire                        merge_ready_o_1_9,

    output      wire        [`DW-1:0]       merge_data_o_1_9,
    output      wire                        merge_valid_o_1_9,
    input       wire                        merge_ready_i_1_9,
    input       wire        [`DW-1:0]       merge_data_i_1_10,
    input       wire                        merge_valid_i_1_10,
    output      wire                        merge_ready_o_1_10,

    output      wire        [`DW-1:0]       merge_data_o_1_10,
    output      wire                        merge_valid_o_1_10,
    input       wire                        merge_ready_i_1_10,
    input       wire        [`DW-1:0]       merge_data_i_1_11,
    input       wire                        merge_valid_i_1_11,
    output      wire                        merge_ready_o_1_11,

    output      wire        [`DW-1:0]       merge_data_o_1_11,
    output      wire                        merge_valid_o_1_11,
    input       wire                        merge_ready_i_1_11,
    input       wire        [`DW-1:0]       merge_data_i_1_12,
    input       wire                        merge_valid_i_1_12,
    output      wire                        merge_ready_o_1_12,

    output      wire        [`DW-1:0]       merge_data_o_1_12,
    output      wire                        merge_valid_o_1_12,
    input       wire                        merge_ready_i_1_12,
    input       wire        [`DW-1:0]       merge_data_i_1_13,
    input       wire                        merge_valid_i_1_13,
    output      wire                        merge_ready_o_1_13,

    output      wire        [`DW-1:0]       merge_data_o_1_13,
    output      wire                        merge_valid_o_1_13,
    input       wire                        merge_ready_i_1_13,
    input       wire        [`DW-1:0]       merge_data_i_1_14,
    input       wire                        merge_valid_i_1_14,
    output      wire                        merge_ready_o_1_14,

    output      wire        [`DW-1:0]       merge_data_o_1_14,
    output      wire                        merge_valid_o_1_14,
    input       wire                        merge_ready_i_1_14,
    input       wire        [`DW-1:0]       merge_data_i_1_15,
    input       wire                        merge_valid_i_1_15,
    output      wire                        merge_ready_o_1_15,

    output      wire        [`DW-1:0]       merge_data_o_1_15,
    output      wire                        merge_valid_o_1_15,
    input       wire                        merge_ready_i_1_15,
    input       wire        [`DW-1:0]       merge_data_i_1_16,
    input       wire                        merge_valid_i_1_16,
    output      wire                        merge_ready_o_1_16,

    output      wire        [`DW-1:0]       merge_data_o_1_16,
    output      wire                        merge_valid_o_1_16,
    input       wire                        merge_ready_i_1_16,
    input       wire        [`DW-1:0]       merge_data_i_1_17,
    input       wire                        merge_valid_i_1_17,
    output      wire                        merge_ready_o_1_17,

    output      wire        [`DW-1:0]       merge_data_o_1_17,
    output      wire                        merge_valid_o_1_17,
    input       wire                        merge_ready_i_1_17,
    input       wire        [`DW-1:0]       merge_data_i_1_18,
    input       wire                        merge_valid_i_1_18,
    output      wire                        merge_ready_o_1_18,

    output      wire        [`DW-1:0]       merge_data_o_1_18,
    output      wire                        merge_valid_o_1_18,
    input       wire                        merge_ready_i_1_18,
    input       wire        [`DW-1:0]       merge_data_i_1_19,
    input       wire                        merge_valid_i_1_19,
    output      wire                        merge_ready_o_1_19,

    output      wire        [`DW-1:0]       merge_data_o_1_19,
    output      wire                        merge_valid_o_1_19,
    input       wire                        merge_ready_i_1_19,
    input       wire        [`DW-1:0]       merge_data_i_1_20,
    input       wire                        merge_valid_i_1_20,
    output      wire                        merge_ready_o_1_20,

    output      wire        [`DW-1:0]       merge_data_o_1_20,
    output      wire                        merge_valid_o_1_20,
    input       wire                        merge_ready_i_1_20,
    input       wire        [`DW-1:0]       merge_data_i_1_21,
    input       wire                        merge_valid_i_1_21,
    output      wire                        merge_ready_o_1_21,

    output      wire        [`DW-1:0]       merge_data_o_1_21,
    output      wire                        merge_valid_o_1_21,
    input       wire                        merge_ready_i_1_21,
    input       wire        [`DW-1:0]       merge_data_i_1_22,
    input       wire                        merge_valid_i_1_22,
    output      wire                        merge_ready_o_1_22,

    output      wire        [`DW-1:0]       merge_data_o_1_22,
    output      wire                        merge_valid_o_1_22,
    input       wire                        merge_ready_i_1_22,
    input       wire        [`DW-1:0]       merge_data_i_1_23,
    input       wire                        merge_valid_i_1_23,
    output      wire                        merge_ready_o_1_23,

    output      wire        [`DW-1:0]       merge_data_o_1_23,
    output      wire                        merge_valid_o_1_23,
    input       wire                        merge_ready_i_1_23,
    input       wire        [`DW-1:0]       merge_data_i_1_24,
    input       wire                        merge_valid_i_1_24,
    output      wire                        merge_ready_o_1_24,

    output      wire        [`DW-1:0]       merge_data_o_1_24,
    output      wire                        merge_valid_o_1_24,
    input       wire                        merge_ready_i_1_24,
    input       wire        [`DW-1:0]       merge_data_i_2_0,
    input       wire                        merge_valid_i_2_0,
    output      wire                        merge_ready_o_2_0,

    output      wire        [`DW-1:0]       merge_data_o_2_0,
    output      wire                        merge_valid_o_2_0,
    input       wire                        merge_ready_i_2_0,
    input       wire        [`DW-1:0]       merge_data_i_2_1,
    input       wire                        merge_valid_i_2_1,
    output      wire                        merge_ready_o_2_1,

    output      wire        [`DW-1:0]       merge_data_o_2_1,
    output      wire                        merge_valid_o_2_1,
    input       wire                        merge_ready_i_2_1,
    input       wire        [`DW-1:0]       merge_data_i_2_2,
    input       wire                        merge_valid_i_2_2,
    output      wire                        merge_ready_o_2_2,

    output      wire        [`DW-1:0]       merge_data_o_2_2,
    output      wire                        merge_valid_o_2_2,
    input       wire                        merge_ready_i_2_2,
    input       wire        [`DW-1:0]       merge_data_i_2_3,
    input       wire                        merge_valid_i_2_3,
    output      wire                        merge_ready_o_2_3,

    output      wire        [`DW-1:0]       merge_data_o_2_3,
    output      wire                        merge_valid_o_2_3,
    input       wire                        merge_ready_i_2_3,
    input       wire        [`DW-1:0]       merge_data_i_2_4,
    input       wire                        merge_valid_i_2_4,
    output      wire                        merge_ready_o_2_4,

    output      wire        [`DW-1:0]       merge_data_o_2_4,
    output      wire                        merge_valid_o_2_4,
    input       wire                        merge_ready_i_2_4,
    input       wire        [`DW-1:0]       merge_data_i_2_5,
    input       wire                        merge_valid_i_2_5,
    output      wire                        merge_ready_o_2_5,

    output      wire        [`DW-1:0]       merge_data_o_2_5,
    output      wire                        merge_valid_o_2_5,
    input       wire                        merge_ready_i_2_5,
    input       wire        [`DW-1:0]       merge_data_i_2_6,
    input       wire                        merge_valid_i_2_6,
    output      wire                        merge_ready_o_2_6,

    output      wire        [`DW-1:0]       merge_data_o_2_6,
    output      wire                        merge_valid_o_2_6,
    input       wire                        merge_ready_i_2_6,
    input       wire        [`DW-1:0]       merge_data_i_2_7,
    input       wire                        merge_valid_i_2_7,
    output      wire                        merge_ready_o_2_7,

    output      wire        [`DW-1:0]       merge_data_o_2_7,
    output      wire                        merge_valid_o_2_7,
    input       wire                        merge_ready_i_2_7,
    input       wire        [`DW-1:0]       merge_data_i_2_8,
    input       wire                        merge_valid_i_2_8,
    output      wire                        merge_ready_o_2_8,

    output      wire        [`DW-1:0]       merge_data_o_2_8,
    output      wire                        merge_valid_o_2_8,
    input       wire                        merge_ready_i_2_8,
    input       wire        [`DW-1:0]       merge_data_i_2_9,
    input       wire                        merge_valid_i_2_9,
    output      wire                        merge_ready_o_2_9,

    output      wire        [`DW-1:0]       merge_data_o_2_9,
    output      wire                        merge_valid_o_2_9,
    input       wire                        merge_ready_i_2_9,
    input       wire        [`DW-1:0]       merge_data_i_2_10,
    input       wire                        merge_valid_i_2_10,
    output      wire                        merge_ready_o_2_10,

    output      wire        [`DW-1:0]       merge_data_o_2_10,
    output      wire                        merge_valid_o_2_10,
    input       wire                        merge_ready_i_2_10,
    input       wire        [`DW-1:0]       merge_data_i_2_11,
    input       wire                        merge_valid_i_2_11,
    output      wire                        merge_ready_o_2_11,

    output      wire        [`DW-1:0]       merge_data_o_2_11,
    output      wire                        merge_valid_o_2_11,
    input       wire                        merge_ready_i_2_11,
    input       wire        [`DW-1:0]       merge_data_i_2_12,
    input       wire                        merge_valid_i_2_12,
    output      wire                        merge_ready_o_2_12,

    output      wire        [`DW-1:0]       merge_data_o_2_12,
    output      wire                        merge_valid_o_2_12,
    input       wire                        merge_ready_i_2_12,
    input       wire        [`DW-1:0]       merge_data_i_2_13,
    input       wire                        merge_valid_i_2_13,
    output      wire                        merge_ready_o_2_13,

    output      wire        [`DW-1:0]       merge_data_o_2_13,
    output      wire                        merge_valid_o_2_13,
    input       wire                        merge_ready_i_2_13,
    input       wire        [`DW-1:0]       merge_data_i_2_14,
    input       wire                        merge_valid_i_2_14,
    output      wire                        merge_ready_o_2_14,

    output      wire        [`DW-1:0]       merge_data_o_2_14,
    output      wire                        merge_valid_o_2_14,
    input       wire                        merge_ready_i_2_14,
    input       wire        [`DW-1:0]       merge_data_i_2_15,
    input       wire                        merge_valid_i_2_15,
    output      wire                        merge_ready_o_2_15,

    output      wire        [`DW-1:0]       merge_data_o_2_15,
    output      wire                        merge_valid_o_2_15,
    input       wire                        merge_ready_i_2_15,
    input       wire        [`DW-1:0]       merge_data_i_2_16,
    input       wire                        merge_valid_i_2_16,
    output      wire                        merge_ready_o_2_16,

    output      wire        [`DW-1:0]       merge_data_o_2_16,
    output      wire                        merge_valid_o_2_16,
    input       wire                        merge_ready_i_2_16,
    input       wire        [`DW-1:0]       merge_data_i_2_17,
    input       wire                        merge_valid_i_2_17,
    output      wire                        merge_ready_o_2_17,

    output      wire        [`DW-1:0]       merge_data_o_2_17,
    output      wire                        merge_valid_o_2_17,
    input       wire                        merge_ready_i_2_17,
    input       wire        [`DW-1:0]       merge_data_i_2_18,
    input       wire                        merge_valid_i_2_18,
    output      wire                        merge_ready_o_2_18,

    output      wire        [`DW-1:0]       merge_data_o_2_18,
    output      wire                        merge_valid_o_2_18,
    input       wire                        merge_ready_i_2_18,
    input       wire        [`DW-1:0]       merge_data_i_2_19,
    input       wire                        merge_valid_i_2_19,
    output      wire                        merge_ready_o_2_19,

    output      wire        [`DW-1:0]       merge_data_o_2_19,
    output      wire                        merge_valid_o_2_19,
    input       wire                        merge_ready_i_2_19,
    input       wire        [`DW-1:0]       merge_data_i_2_20,
    input       wire                        merge_valid_i_2_20,
    output      wire                        merge_ready_o_2_20,

    output      wire        [`DW-1:0]       merge_data_o_2_20,
    output      wire                        merge_valid_o_2_20,
    input       wire                        merge_ready_i_2_20,
    input       wire        [`DW-1:0]       merge_data_i_2_21,
    input       wire                        merge_valid_i_2_21,
    output      wire                        merge_ready_o_2_21,

    output      wire        [`DW-1:0]       merge_data_o_2_21,
    output      wire                        merge_valid_o_2_21,
    input       wire                        merge_ready_i_2_21,
    input       wire        [`DW-1:0]       merge_data_i_2_22,
    input       wire                        merge_valid_i_2_22,
    output      wire                        merge_ready_o_2_22,

    output      wire        [`DW-1:0]       merge_data_o_2_22,
    output      wire                        merge_valid_o_2_22,
    input       wire                        merge_ready_i_2_22,
    input       wire        [`DW-1:0]       merge_data_i_2_23,
    input       wire                        merge_valid_i_2_23,
    output      wire                        merge_ready_o_2_23,

    output      wire        [`DW-1:0]       merge_data_o_2_23,
    output      wire                        merge_valid_o_2_23,
    input       wire                        merge_ready_i_2_23,
    input       wire        [`DW-1:0]       merge_data_i_2_24,
    input       wire                        merge_valid_i_2_24,
    output      wire                        merge_ready_o_2_24,

    output      wire        [`DW-1:0]       merge_data_o_2_24,
    output      wire                        merge_valid_o_2_24,
    input       wire                        merge_ready_i_2_24,
    input       wire        [`DW-1:0]       merge_data_i_3_0,
    input       wire                        merge_valid_i_3_0,
    output      wire                        merge_ready_o_3_0,

    output      wire        [`DW-1:0]       merge_data_o_3_0,
    output      wire                        merge_valid_o_3_0,
    input       wire                        merge_ready_i_3_0,
    input       wire        [`DW-1:0]       merge_data_i_3_1,
    input       wire                        merge_valid_i_3_1,
    output      wire                        merge_ready_o_3_1,

    output      wire        [`DW-1:0]       merge_data_o_3_1,
    output      wire                        merge_valid_o_3_1,
    input       wire                        merge_ready_i_3_1,
    input       wire        [`DW-1:0]       merge_data_i_3_2,
    input       wire                        merge_valid_i_3_2,
    output      wire                        merge_ready_o_3_2,

    output      wire        [`DW-1:0]       merge_data_o_3_2,
    output      wire                        merge_valid_o_3_2,
    input       wire                        merge_ready_i_3_2,
    input       wire        [`DW-1:0]       merge_data_i_3_3,
    input       wire                        merge_valid_i_3_3,
    output      wire                        merge_ready_o_3_3,

    output      wire        [`DW-1:0]       merge_data_o_3_3,
    output      wire                        merge_valid_o_3_3,
    input       wire                        merge_ready_i_3_3,
    input       wire        [`DW-1:0]       merge_data_i_3_4,
    input       wire                        merge_valid_i_3_4,
    output      wire                        merge_ready_o_3_4,

    output      wire        [`DW-1:0]       merge_data_o_3_4,
    output      wire                        merge_valid_o_3_4,
    input       wire                        merge_ready_i_3_4,
    input       wire        [`DW-1:0]       merge_data_i_3_5,
    input       wire                        merge_valid_i_3_5,
    output      wire                        merge_ready_o_3_5,

    output      wire        [`DW-1:0]       merge_data_o_3_5,
    output      wire                        merge_valid_o_3_5,
    input       wire                        merge_ready_i_3_5,
    input       wire        [`DW-1:0]       merge_data_i_3_6,
    input       wire                        merge_valid_i_3_6,
    output      wire                        merge_ready_o_3_6,

    output      wire        [`DW-1:0]       merge_data_o_3_6,
    output      wire                        merge_valid_o_3_6,
    input       wire                        merge_ready_i_3_6,
    input       wire        [`DW-1:0]       merge_data_i_3_7,
    input       wire                        merge_valid_i_3_7,
    output      wire                        merge_ready_o_3_7,

    output      wire        [`DW-1:0]       merge_data_o_3_7,
    output      wire                        merge_valid_o_3_7,
    input       wire                        merge_ready_i_3_7,
    input       wire        [`DW-1:0]       merge_data_i_3_8,
    input       wire                        merge_valid_i_3_8,
    output      wire                        merge_ready_o_3_8,

    output      wire        [`DW-1:0]       merge_data_o_3_8,
    output      wire                        merge_valid_o_3_8,
    input       wire                        merge_ready_i_3_8,
    input       wire        [`DW-1:0]       merge_data_i_3_9,
    input       wire                        merge_valid_i_3_9,
    output      wire                        merge_ready_o_3_9,

    output      wire        [`DW-1:0]       merge_data_o_3_9,
    output      wire                        merge_valid_o_3_9,
    input       wire                        merge_ready_i_3_9,
    input       wire        [`DW-1:0]       merge_data_i_3_10,
    input       wire                        merge_valid_i_3_10,
    output      wire                        merge_ready_o_3_10,

    output      wire        [`DW-1:0]       merge_data_o_3_10,
    output      wire                        merge_valid_o_3_10,
    input       wire                        merge_ready_i_3_10,
    input       wire        [`DW-1:0]       merge_data_i_3_11,
    input       wire                        merge_valid_i_3_11,
    output      wire                        merge_ready_o_3_11,

    output      wire        [`DW-1:0]       merge_data_o_3_11,
    output      wire                        merge_valid_o_3_11,
    input       wire                        merge_ready_i_3_11,
    input       wire        [`DW-1:0]       merge_data_i_3_12,
    input       wire                        merge_valid_i_3_12,
    output      wire                        merge_ready_o_3_12,

    output      wire        [`DW-1:0]       merge_data_o_3_12,
    output      wire                        merge_valid_o_3_12,
    input       wire                        merge_ready_i_3_12,
    input       wire        [`DW-1:0]       merge_data_i_3_13,
    input       wire                        merge_valid_i_3_13,
    output      wire                        merge_ready_o_3_13,

    output      wire        [`DW-1:0]       merge_data_o_3_13,
    output      wire                        merge_valid_o_3_13,
    input       wire                        merge_ready_i_3_13,
    input       wire        [`DW-1:0]       merge_data_i_3_14,
    input       wire                        merge_valid_i_3_14,
    output      wire                        merge_ready_o_3_14,

    output      wire        [`DW-1:0]       merge_data_o_3_14,
    output      wire                        merge_valid_o_3_14,
    input       wire                        merge_ready_i_3_14,
    input       wire        [`DW-1:0]       merge_data_i_3_15,
    input       wire                        merge_valid_i_3_15,
    output      wire                        merge_ready_o_3_15,

    output      wire        [`DW-1:0]       merge_data_o_3_15,
    output      wire                        merge_valid_o_3_15,
    input       wire                        merge_ready_i_3_15,
    input       wire        [`DW-1:0]       merge_data_i_3_16,
    input       wire                        merge_valid_i_3_16,
    output      wire                        merge_ready_o_3_16,

    output      wire        [`DW-1:0]       merge_data_o_3_16,
    output      wire                        merge_valid_o_3_16,
    input       wire                        merge_ready_i_3_16,
    input       wire        [`DW-1:0]       merge_data_i_3_17,
    input       wire                        merge_valid_i_3_17,
    output      wire                        merge_ready_o_3_17,

    output      wire        [`DW-1:0]       merge_data_o_3_17,
    output      wire                        merge_valid_o_3_17,
    input       wire                        merge_ready_i_3_17,
    input       wire        [`DW-1:0]       merge_data_i_3_18,
    input       wire                        merge_valid_i_3_18,
    output      wire                        merge_ready_o_3_18,

    output      wire        [`DW-1:0]       merge_data_o_3_18,
    output      wire                        merge_valid_o_3_18,
    input       wire                        merge_ready_i_3_18,
    input       wire        [`DW-1:0]       merge_data_i_3_19,
    input       wire                        merge_valid_i_3_19,
    output      wire                        merge_ready_o_3_19,

    output      wire        [`DW-1:0]       merge_data_o_3_19,
    output      wire                        merge_valid_o_3_19,
    input       wire                        merge_ready_i_3_19,
    input       wire        [`DW-1:0]       merge_data_i_3_20,
    input       wire                        merge_valid_i_3_20,
    output      wire                        merge_ready_o_3_20,

    output      wire        [`DW-1:0]       merge_data_o_3_20,
    output      wire                        merge_valid_o_3_20,
    input       wire                        merge_ready_i_3_20,
    input       wire        [`DW-1:0]       merge_data_i_3_21,
    input       wire                        merge_valid_i_3_21,
    output      wire                        merge_ready_o_3_21,

    output      wire        [`DW-1:0]       merge_data_o_3_21,
    output      wire                        merge_valid_o_3_21,
    input       wire                        merge_ready_i_3_21,
    input       wire        [`DW-1:0]       merge_data_i_3_22,
    input       wire                        merge_valid_i_3_22,
    output      wire                        merge_ready_o_3_22,

    output      wire        [`DW-1:0]       merge_data_o_3_22,
    output      wire                        merge_valid_o_3_22,
    input       wire                        merge_ready_i_3_22,
    input       wire        [`DW-1:0]       merge_data_i_3_23,
    input       wire                        merge_valid_i_3_23,
    output      wire                        merge_ready_o_3_23,

    output      wire        [`DW-1:0]       merge_data_o_3_23,
    output      wire                        merge_valid_o_3_23,
    input       wire                        merge_ready_i_3_23,
    input       wire        [`DW-1:0]       merge_data_i_3_24,
    input       wire                        merge_valid_i_3_24,
    output      wire                        merge_ready_o_3_24,

    output      wire        [`DW-1:0]       merge_data_o_3_24,
    output      wire                        merge_valid_o_3_24,
    input       wire                        merge_ready_i_3_24,
    input       wire        [`DW-1:0]       merge_data_i_4_0,
    input       wire                        merge_valid_i_4_0,
    output      wire                        merge_ready_o_4_0,

    output      wire        [`DW-1:0]       merge_data_o_4_0,
    output      wire                        merge_valid_o_4_0,
    input       wire                        merge_ready_i_4_0,
    input       wire        [`DW-1:0]       merge_data_i_4_1,
    input       wire                        merge_valid_i_4_1,
    output      wire                        merge_ready_o_4_1,

    output      wire        [`DW-1:0]       merge_data_o_4_1,
    output      wire                        merge_valid_o_4_1,
    input       wire                        merge_ready_i_4_1,
    input       wire        [`DW-1:0]       merge_data_i_4_2,
    input       wire                        merge_valid_i_4_2,
    output      wire                        merge_ready_o_4_2,

    output      wire        [`DW-1:0]       merge_data_o_4_2,
    output      wire                        merge_valid_o_4_2,
    input       wire                        merge_ready_i_4_2,
    input       wire        [`DW-1:0]       merge_data_i_4_3,
    input       wire                        merge_valid_i_4_3,
    output      wire                        merge_ready_o_4_3,

    output      wire        [`DW-1:0]       merge_data_o_4_3,
    output      wire                        merge_valid_o_4_3,
    input       wire                        merge_ready_i_4_3,
    input       wire        [`DW-1:0]       merge_data_i_4_4,
    input       wire                        merge_valid_i_4_4,
    output      wire                        merge_ready_o_4_4,

    output      wire        [`DW-1:0]       merge_data_o_4_4,
    output      wire                        merge_valid_o_4_4,
    input       wire                        merge_ready_i_4_4,
    input       wire        [`DW-1:0]       merge_data_i_4_5,
    input       wire                        merge_valid_i_4_5,
    output      wire                        merge_ready_o_4_5,

    output      wire        [`DW-1:0]       merge_data_o_4_5,
    output      wire                        merge_valid_o_4_5,
    input       wire                        merge_ready_i_4_5,
    input       wire        [`DW-1:0]       merge_data_i_4_6,
    input       wire                        merge_valid_i_4_6,
    output      wire                        merge_ready_o_4_6,

    output      wire        [`DW-1:0]       merge_data_o_4_6,
    output      wire                        merge_valid_o_4_6,
    input       wire                        merge_ready_i_4_6,
    input       wire        [`DW-1:0]       merge_data_i_4_7,
    input       wire                        merge_valid_i_4_7,
    output      wire                        merge_ready_o_4_7,

    output      wire        [`DW-1:0]       merge_data_o_4_7,
    output      wire                        merge_valid_o_4_7,
    input       wire                        merge_ready_i_4_7,
    input       wire        [`DW-1:0]       merge_data_i_4_8,
    input       wire                        merge_valid_i_4_8,
    output      wire                        merge_ready_o_4_8,

    output      wire        [`DW-1:0]       merge_data_o_4_8,
    output      wire                        merge_valid_o_4_8,
    input       wire                        merge_ready_i_4_8,
    input       wire        [`DW-1:0]       merge_data_i_4_9,
    input       wire                        merge_valid_i_4_9,
    output      wire                        merge_ready_o_4_9,

    output      wire        [`DW-1:0]       merge_data_o_4_9,
    output      wire                        merge_valid_o_4_9,
    input       wire                        merge_ready_i_4_9,
    input       wire        [`DW-1:0]       merge_data_i_4_10,
    input       wire                        merge_valid_i_4_10,
    output      wire                        merge_ready_o_4_10,

    output      wire        [`DW-1:0]       merge_data_o_4_10,
    output      wire                        merge_valid_o_4_10,
    input       wire                        merge_ready_i_4_10,
    input       wire        [`DW-1:0]       merge_data_i_4_11,
    input       wire                        merge_valid_i_4_11,
    output      wire                        merge_ready_o_4_11,

    output      wire        [`DW-1:0]       merge_data_o_4_11,
    output      wire                        merge_valid_o_4_11,
    input       wire                        merge_ready_i_4_11,
    input       wire        [`DW-1:0]       merge_data_i_4_12,
    input       wire                        merge_valid_i_4_12,
    output      wire                        merge_ready_o_4_12,

    output      wire        [`DW-1:0]       merge_data_o_4_12,
    output      wire                        merge_valid_o_4_12,
    input       wire                        merge_ready_i_4_12,
    input       wire        [`DW-1:0]       merge_data_i_4_13,
    input       wire                        merge_valid_i_4_13,
    output      wire                        merge_ready_o_4_13,

    output      wire        [`DW-1:0]       merge_data_o_4_13,
    output      wire                        merge_valid_o_4_13,
    input       wire                        merge_ready_i_4_13,
    input       wire        [`DW-1:0]       merge_data_i_4_14,
    input       wire                        merge_valid_i_4_14,
    output      wire                        merge_ready_o_4_14,

    output      wire        [`DW-1:0]       merge_data_o_4_14,
    output      wire                        merge_valid_o_4_14,
    input       wire                        merge_ready_i_4_14,
    input       wire        [`DW-1:0]       merge_data_i_4_15,
    input       wire                        merge_valid_i_4_15,
    output      wire                        merge_ready_o_4_15,

    output      wire        [`DW-1:0]       merge_data_o_4_15,
    output      wire                        merge_valid_o_4_15,
    input       wire                        merge_ready_i_4_15,
    input       wire        [`DW-1:0]       merge_data_i_4_16,
    input       wire                        merge_valid_i_4_16,
    output      wire                        merge_ready_o_4_16,

    output      wire        [`DW-1:0]       merge_data_o_4_16,
    output      wire                        merge_valid_o_4_16,
    input       wire                        merge_ready_i_4_16,
    input       wire        [`DW-1:0]       merge_data_i_4_17,
    input       wire                        merge_valid_i_4_17,
    output      wire                        merge_ready_o_4_17,

    output      wire        [`DW-1:0]       merge_data_o_4_17,
    output      wire                        merge_valid_o_4_17,
    input       wire                        merge_ready_i_4_17,
    input       wire        [`DW-1:0]       merge_data_i_4_18,
    input       wire                        merge_valid_i_4_18,
    output      wire                        merge_ready_o_4_18,

    output      wire        [`DW-1:0]       merge_data_o_4_18,
    output      wire                        merge_valid_o_4_18,
    input       wire                        merge_ready_i_4_18,
    input       wire        [`DW-1:0]       merge_data_i_4_19,
    input       wire                        merge_valid_i_4_19,
    output      wire                        merge_ready_o_4_19,

    output      wire        [`DW-1:0]       merge_data_o_4_19,
    output      wire                        merge_valid_o_4_19,
    input       wire                        merge_ready_i_4_19,
    input       wire        [`DW-1:0]       merge_data_i_4_20,
    input       wire                        merge_valid_i_4_20,
    output      wire                        merge_ready_o_4_20,

    output      wire        [`DW-1:0]       merge_data_o_4_20,
    output      wire                        merge_valid_o_4_20,
    input       wire                        merge_ready_i_4_20,
    input       wire        [`DW-1:0]       merge_data_i_4_21,
    input       wire                        merge_valid_i_4_21,
    output      wire                        merge_ready_o_4_21,

    output      wire        [`DW-1:0]       merge_data_o_4_21,
    output      wire                        merge_valid_o_4_21,
    input       wire                        merge_ready_i_4_21,
    input       wire        [`DW-1:0]       merge_data_i_4_22,
    input       wire                        merge_valid_i_4_22,
    output      wire                        merge_ready_o_4_22,

    output      wire        [`DW-1:0]       merge_data_o_4_22,
    output      wire                        merge_valid_o_4_22,
    input       wire                        merge_ready_i_4_22,
    input       wire        [`DW-1:0]       merge_data_i_4_23,
    input       wire                        merge_valid_i_4_23,
    output      wire                        merge_ready_o_4_23,

    output      wire        [`DW-1:0]       merge_data_o_4_23,
    output      wire                        merge_valid_o_4_23,
    input       wire                        merge_ready_i_4_23,
    input       wire        [`DW-1:0]       merge_data_i_4_24,
    input       wire                        merge_valid_i_4_24,
    output      wire                        merge_ready_o_4_24,

    output      wire        [`DW-1:0]       merge_data_o_4_24,
    output      wire                        merge_valid_o_4_24,
    input       wire                        merge_ready_i_4_24,
    input       wire        [`DW-1:0]       merge_data_i_5_0,
    input       wire                        merge_valid_i_5_0,
    output      wire                        merge_ready_o_5_0,

    output      wire        [`DW-1:0]       merge_data_o_5_0,
    output      wire                        merge_valid_o_5_0,
    input       wire                        merge_ready_i_5_0,
    input       wire        [`DW-1:0]       merge_data_i_5_1,
    input       wire                        merge_valid_i_5_1,
    output      wire                        merge_ready_o_5_1,

    output      wire        [`DW-1:0]       merge_data_o_5_1,
    output      wire                        merge_valid_o_5_1,
    input       wire                        merge_ready_i_5_1,
    input       wire        [`DW-1:0]       merge_data_i_5_2,
    input       wire                        merge_valid_i_5_2,
    output      wire                        merge_ready_o_5_2,

    output      wire        [`DW-1:0]       merge_data_o_5_2,
    output      wire                        merge_valid_o_5_2,
    input       wire                        merge_ready_i_5_2,
    input       wire        [`DW-1:0]       merge_data_i_5_3,
    input       wire                        merge_valid_i_5_3,
    output      wire                        merge_ready_o_5_3,

    output      wire        [`DW-1:0]       merge_data_o_5_3,
    output      wire                        merge_valid_o_5_3,
    input       wire                        merge_ready_i_5_3,
    input       wire        [`DW-1:0]       merge_data_i_5_4,
    input       wire                        merge_valid_i_5_4,
    output      wire                        merge_ready_o_5_4,

    output      wire        [`DW-1:0]       merge_data_o_5_4,
    output      wire                        merge_valid_o_5_4,
    input       wire                        merge_ready_i_5_4,
    input       wire        [`DW-1:0]       merge_data_i_5_5,
    input       wire                        merge_valid_i_5_5,
    output      wire                        merge_ready_o_5_5,

    output      wire        [`DW-1:0]       merge_data_o_5_5,
    output      wire                        merge_valid_o_5_5,
    input       wire                        merge_ready_i_5_5,
    input       wire        [`DW-1:0]       merge_data_i_5_6,
    input       wire                        merge_valid_i_5_6,
    output      wire                        merge_ready_o_5_6,

    output      wire        [`DW-1:0]       merge_data_o_5_6,
    output      wire                        merge_valid_o_5_6,
    input       wire                        merge_ready_i_5_6,
    input       wire        [`DW-1:0]       merge_data_i_5_7,
    input       wire                        merge_valid_i_5_7,
    output      wire                        merge_ready_o_5_7,

    output      wire        [`DW-1:0]       merge_data_o_5_7,
    output      wire                        merge_valid_o_5_7,
    input       wire                        merge_ready_i_5_7,
    input       wire        [`DW-1:0]       merge_data_i_5_8,
    input       wire                        merge_valid_i_5_8,
    output      wire                        merge_ready_o_5_8,

    output      wire        [`DW-1:0]       merge_data_o_5_8,
    output      wire                        merge_valid_o_5_8,
    input       wire                        merge_ready_i_5_8,
    input       wire        [`DW-1:0]       merge_data_i_5_9,
    input       wire                        merge_valid_i_5_9,
    output      wire                        merge_ready_o_5_9,

    output      wire        [`DW-1:0]       merge_data_o_5_9,
    output      wire                        merge_valid_o_5_9,
    input       wire                        merge_ready_i_5_9,
    input       wire        [`DW-1:0]       merge_data_i_5_10,
    input       wire                        merge_valid_i_5_10,
    output      wire                        merge_ready_o_5_10,

    output      wire        [`DW-1:0]       merge_data_o_5_10,
    output      wire                        merge_valid_o_5_10,
    input       wire                        merge_ready_i_5_10,
    input       wire        [`DW-1:0]       merge_data_i_5_11,
    input       wire                        merge_valid_i_5_11,
    output      wire                        merge_ready_o_5_11,

    output      wire        [`DW-1:0]       merge_data_o_5_11,
    output      wire                        merge_valid_o_5_11,
    input       wire                        merge_ready_i_5_11,
    input       wire        [`DW-1:0]       merge_data_i_5_12,
    input       wire                        merge_valid_i_5_12,
    output      wire                        merge_ready_o_5_12,

    output      wire        [`DW-1:0]       merge_data_o_5_12,
    output      wire                        merge_valid_o_5_12,
    input       wire                        merge_ready_i_5_12,
    input       wire        [`DW-1:0]       merge_data_i_5_13,
    input       wire                        merge_valid_i_5_13,
    output      wire                        merge_ready_o_5_13,

    output      wire        [`DW-1:0]       merge_data_o_5_13,
    output      wire                        merge_valid_o_5_13,
    input       wire                        merge_ready_i_5_13,
    input       wire        [`DW-1:0]       merge_data_i_5_14,
    input       wire                        merge_valid_i_5_14,
    output      wire                        merge_ready_o_5_14,

    output      wire        [`DW-1:0]       merge_data_o_5_14,
    output      wire                        merge_valid_o_5_14,
    input       wire                        merge_ready_i_5_14,
    input       wire        [`DW-1:0]       merge_data_i_5_15,
    input       wire                        merge_valid_i_5_15,
    output      wire                        merge_ready_o_5_15,

    output      wire        [`DW-1:0]       merge_data_o_5_15,
    output      wire                        merge_valid_o_5_15,
    input       wire                        merge_ready_i_5_15,
    input       wire        [`DW-1:0]       merge_data_i_5_16,
    input       wire                        merge_valid_i_5_16,
    output      wire                        merge_ready_o_5_16,

    output      wire        [`DW-1:0]       merge_data_o_5_16,
    output      wire                        merge_valid_o_5_16,
    input       wire                        merge_ready_i_5_16,
    input       wire        [`DW-1:0]       merge_data_i_5_17,
    input       wire                        merge_valid_i_5_17,
    output      wire                        merge_ready_o_5_17,

    output      wire        [`DW-1:0]       merge_data_o_5_17,
    output      wire                        merge_valid_o_5_17,
    input       wire                        merge_ready_i_5_17,
    input       wire        [`DW-1:0]       merge_data_i_5_18,
    input       wire                        merge_valid_i_5_18,
    output      wire                        merge_ready_o_5_18,

    output      wire        [`DW-1:0]       merge_data_o_5_18,
    output      wire                        merge_valid_o_5_18,
    input       wire                        merge_ready_i_5_18,
    input       wire        [`DW-1:0]       merge_data_i_5_19,
    input       wire                        merge_valid_i_5_19,
    output      wire                        merge_ready_o_5_19,

    output      wire        [`DW-1:0]       merge_data_o_5_19,
    output      wire                        merge_valid_o_5_19,
    input       wire                        merge_ready_i_5_19,
    input       wire        [`DW-1:0]       merge_data_i_5_20,
    input       wire                        merge_valid_i_5_20,
    output      wire                        merge_ready_o_5_20,

    output      wire        [`DW-1:0]       merge_data_o_5_20,
    output      wire                        merge_valid_o_5_20,
    input       wire                        merge_ready_i_5_20,
    input       wire        [`DW-1:0]       merge_data_i_5_21,
    input       wire                        merge_valid_i_5_21,
    output      wire                        merge_ready_o_5_21,

    output      wire        [`DW-1:0]       merge_data_o_5_21,
    output      wire                        merge_valid_o_5_21,
    input       wire                        merge_ready_i_5_21,
    input       wire        [`DW-1:0]       merge_data_i_5_22,
    input       wire                        merge_valid_i_5_22,
    output      wire                        merge_ready_o_5_22,

    output      wire        [`DW-1:0]       merge_data_o_5_22,
    output      wire                        merge_valid_o_5_22,
    input       wire                        merge_ready_i_5_22,
    input       wire        [`DW-1:0]       merge_data_i_5_23,
    input       wire                        merge_valid_i_5_23,
    output      wire                        merge_ready_o_5_23,

    output      wire        [`DW-1:0]       merge_data_o_5_23,
    output      wire                        merge_valid_o_5_23,
    input       wire                        merge_ready_i_5_23,
    input       wire        [`DW-1:0]       merge_data_i_5_24,
    input       wire                        merge_valid_i_5_24,
    output      wire                        merge_ready_o_5_24,

    output      wire        [`DW-1:0]       merge_data_o_5_24,
    output      wire                        merge_valid_o_5_24,
    input       wire                        merge_ready_i_5_24,
    input       wire        [`DW-1:0]       merge_data_i_6_0,
    input       wire                        merge_valid_i_6_0,
    output      wire                        merge_ready_o_6_0,

    output      wire        [`DW-1:0]       merge_data_o_6_0,
    output      wire                        merge_valid_o_6_0,
    input       wire                        merge_ready_i_6_0,
    input       wire        [`DW-1:0]       merge_data_i_6_1,
    input       wire                        merge_valid_i_6_1,
    output      wire                        merge_ready_o_6_1,

    output      wire        [`DW-1:0]       merge_data_o_6_1,
    output      wire                        merge_valid_o_6_1,
    input       wire                        merge_ready_i_6_1,
    input       wire        [`DW-1:0]       merge_data_i_6_2,
    input       wire                        merge_valid_i_6_2,
    output      wire                        merge_ready_o_6_2,

    output      wire        [`DW-1:0]       merge_data_o_6_2,
    output      wire                        merge_valid_o_6_2,
    input       wire                        merge_ready_i_6_2,
    input       wire        [`DW-1:0]       merge_data_i_6_3,
    input       wire                        merge_valid_i_6_3,
    output      wire                        merge_ready_o_6_3,

    output      wire        [`DW-1:0]       merge_data_o_6_3,
    output      wire                        merge_valid_o_6_3,
    input       wire                        merge_ready_i_6_3,
    input       wire        [`DW-1:0]       merge_data_i_6_4,
    input       wire                        merge_valid_i_6_4,
    output      wire                        merge_ready_o_6_4,

    output      wire        [`DW-1:0]       merge_data_o_6_4,
    output      wire                        merge_valid_o_6_4,
    input       wire                        merge_ready_i_6_4,
    input       wire        [`DW-1:0]       merge_data_i_6_5,
    input       wire                        merge_valid_i_6_5,
    output      wire                        merge_ready_o_6_5,

    output      wire        [`DW-1:0]       merge_data_o_6_5,
    output      wire                        merge_valid_o_6_5,
    input       wire                        merge_ready_i_6_5,
    input       wire        [`DW-1:0]       merge_data_i_6_6,
    input       wire                        merge_valid_i_6_6,
    output      wire                        merge_ready_o_6_6,

    output      wire        [`DW-1:0]       merge_data_o_6_6,
    output      wire                        merge_valid_o_6_6,
    input       wire                        merge_ready_i_6_6,
    input       wire        [`DW-1:0]       merge_data_i_6_7,
    input       wire                        merge_valid_i_6_7,
    output      wire                        merge_ready_o_6_7,

    output      wire        [`DW-1:0]       merge_data_o_6_7,
    output      wire                        merge_valid_o_6_7,
    input       wire                        merge_ready_i_6_7,
    input       wire        [`DW-1:0]       merge_data_i_6_8,
    input       wire                        merge_valid_i_6_8,
    output      wire                        merge_ready_o_6_8,

    output      wire        [`DW-1:0]       merge_data_o_6_8,
    output      wire                        merge_valid_o_6_8,
    input       wire                        merge_ready_i_6_8,
    input       wire        [`DW-1:0]       merge_data_i_6_9,
    input       wire                        merge_valid_i_6_9,
    output      wire                        merge_ready_o_6_9,

    output      wire        [`DW-1:0]       merge_data_o_6_9,
    output      wire                        merge_valid_o_6_9,
    input       wire                        merge_ready_i_6_9,
    input       wire        [`DW-1:0]       merge_data_i_6_10,
    input       wire                        merge_valid_i_6_10,
    output      wire                        merge_ready_o_6_10,

    output      wire        [`DW-1:0]       merge_data_o_6_10,
    output      wire                        merge_valid_o_6_10,
    input       wire                        merge_ready_i_6_10,
    input       wire        [`DW-1:0]       merge_data_i_6_11,
    input       wire                        merge_valid_i_6_11,
    output      wire                        merge_ready_o_6_11,

    output      wire        [`DW-1:0]       merge_data_o_6_11,
    output      wire                        merge_valid_o_6_11,
    input       wire                        merge_ready_i_6_11,
    input       wire        [`DW-1:0]       merge_data_i_6_12,
    input       wire                        merge_valid_i_6_12,
    output      wire                        merge_ready_o_6_12,

    output      wire        [`DW-1:0]       merge_data_o_6_12,
    output      wire                        merge_valid_o_6_12,
    input       wire                        merge_ready_i_6_12,
    input       wire        [`DW-1:0]       merge_data_i_6_13,
    input       wire                        merge_valid_i_6_13,
    output      wire                        merge_ready_o_6_13,

    output      wire        [`DW-1:0]       merge_data_o_6_13,
    output      wire                        merge_valid_o_6_13,
    input       wire                        merge_ready_i_6_13,
    input       wire        [`DW-1:0]       merge_data_i_6_14,
    input       wire                        merge_valid_i_6_14,
    output      wire                        merge_ready_o_6_14,

    output      wire        [`DW-1:0]       merge_data_o_6_14,
    output      wire                        merge_valid_o_6_14,
    input       wire                        merge_ready_i_6_14,
    input       wire        [`DW-1:0]       merge_data_i_6_15,
    input       wire                        merge_valid_i_6_15,
    output      wire                        merge_ready_o_6_15,

    output      wire        [`DW-1:0]       merge_data_o_6_15,
    output      wire                        merge_valid_o_6_15,
    input       wire                        merge_ready_i_6_15,
    input       wire        [`DW-1:0]       merge_data_i_6_16,
    input       wire                        merge_valid_i_6_16,
    output      wire                        merge_ready_o_6_16,

    output      wire        [`DW-1:0]       merge_data_o_6_16,
    output      wire                        merge_valid_o_6_16,
    input       wire                        merge_ready_i_6_16,
    input       wire        [`DW-1:0]       merge_data_i_6_17,
    input       wire                        merge_valid_i_6_17,
    output      wire                        merge_ready_o_6_17,

    output      wire        [`DW-1:0]       merge_data_o_6_17,
    output      wire                        merge_valid_o_6_17,
    input       wire                        merge_ready_i_6_17,
    input       wire        [`DW-1:0]       merge_data_i_6_18,
    input       wire                        merge_valid_i_6_18,
    output      wire                        merge_ready_o_6_18,

    output      wire        [`DW-1:0]       merge_data_o_6_18,
    output      wire                        merge_valid_o_6_18,
    input       wire                        merge_ready_i_6_18,
    input       wire        [`DW-1:0]       merge_data_i_6_19,
    input       wire                        merge_valid_i_6_19,
    output      wire                        merge_ready_o_6_19,

    output      wire        [`DW-1:0]       merge_data_o_6_19,
    output      wire                        merge_valid_o_6_19,
    input       wire                        merge_ready_i_6_19,
    input       wire        [`DW-1:0]       merge_data_i_6_20,
    input       wire                        merge_valid_i_6_20,
    output      wire                        merge_ready_o_6_20,

    output      wire        [`DW-1:0]       merge_data_o_6_20,
    output      wire                        merge_valid_o_6_20,
    input       wire                        merge_ready_i_6_20,
    input       wire        [`DW-1:0]       merge_data_i_6_21,
    input       wire                        merge_valid_i_6_21,
    output      wire                        merge_ready_o_6_21,

    output      wire        [`DW-1:0]       merge_data_o_6_21,
    output      wire                        merge_valid_o_6_21,
    input       wire                        merge_ready_i_6_21,
    input       wire        [`DW-1:0]       merge_data_i_6_22,
    input       wire                        merge_valid_i_6_22,
    output      wire                        merge_ready_o_6_22,

    output      wire        [`DW-1:0]       merge_data_o_6_22,
    output      wire                        merge_valid_o_6_22,
    input       wire                        merge_ready_i_6_22,
    input       wire        [`DW-1:0]       merge_data_i_6_23,
    input       wire                        merge_valid_i_6_23,
    output      wire                        merge_ready_o_6_23,

    output      wire        [`DW-1:0]       merge_data_o_6_23,
    output      wire                        merge_valid_o_6_23,
    input       wire                        merge_ready_i_6_23,
    input       wire        [`DW-1:0]       merge_data_i_6_24,
    input       wire                        merge_valid_i_6_24,
    output      wire                        merge_ready_o_6_24,

    output      wire        [`DW-1:0]       merge_data_o_6_24,
    output      wire                        merge_valid_o_6_24,
    input       wire                        merge_ready_i_6_24,
    input       wire        [`DW-1:0]       merge_data_i_7_0,
    input       wire                        merge_valid_i_7_0,
    output      wire                        merge_ready_o_7_0,

    output      wire        [`DW-1:0]       merge_data_o_7_0,
    output      wire                        merge_valid_o_7_0,
    input       wire                        merge_ready_i_7_0,
    input       wire        [`DW-1:0]       merge_data_i_7_1,
    input       wire                        merge_valid_i_7_1,
    output      wire                        merge_ready_o_7_1,

    output      wire        [`DW-1:0]       merge_data_o_7_1,
    output      wire                        merge_valid_o_7_1,
    input       wire                        merge_ready_i_7_1,
    input       wire        [`DW-1:0]       merge_data_i_7_2,
    input       wire                        merge_valid_i_7_2,
    output      wire                        merge_ready_o_7_2,

    output      wire        [`DW-1:0]       merge_data_o_7_2,
    output      wire                        merge_valid_o_7_2,
    input       wire                        merge_ready_i_7_2,
    input       wire        [`DW-1:0]       merge_data_i_7_3,
    input       wire                        merge_valid_i_7_3,
    output      wire                        merge_ready_o_7_3,

    output      wire        [`DW-1:0]       merge_data_o_7_3,
    output      wire                        merge_valid_o_7_3,
    input       wire                        merge_ready_i_7_3,
    input       wire        [`DW-1:0]       merge_data_i_7_4,
    input       wire                        merge_valid_i_7_4,
    output      wire                        merge_ready_o_7_4,

    output      wire        [`DW-1:0]       merge_data_o_7_4,
    output      wire                        merge_valid_o_7_4,
    input       wire                        merge_ready_i_7_4,
    input       wire        [`DW-1:0]       merge_data_i_7_5,
    input       wire                        merge_valid_i_7_5,
    output      wire                        merge_ready_o_7_5,

    output      wire        [`DW-1:0]       merge_data_o_7_5,
    output      wire                        merge_valid_o_7_5,
    input       wire                        merge_ready_i_7_5,
    input       wire        [`DW-1:0]       merge_data_i_7_6,
    input       wire                        merge_valid_i_7_6,
    output      wire                        merge_ready_o_7_6,

    output      wire        [`DW-1:0]       merge_data_o_7_6,
    output      wire                        merge_valid_o_7_6,
    input       wire                        merge_ready_i_7_6,
    input       wire        [`DW-1:0]       merge_data_i_7_7,
    input       wire                        merge_valid_i_7_7,
    output      wire                        merge_ready_o_7_7,

    output      wire        [`DW-1:0]       merge_data_o_7_7,
    output      wire                        merge_valid_o_7_7,
    input       wire                        merge_ready_i_7_7,
    input       wire        [`DW-1:0]       merge_data_i_7_8,
    input       wire                        merge_valid_i_7_8,
    output      wire                        merge_ready_o_7_8,

    output      wire        [`DW-1:0]       merge_data_o_7_8,
    output      wire                        merge_valid_o_7_8,
    input       wire                        merge_ready_i_7_8,
    input       wire        [`DW-1:0]       merge_data_i_7_9,
    input       wire                        merge_valid_i_7_9,
    output      wire                        merge_ready_o_7_9,

    output      wire        [`DW-1:0]       merge_data_o_7_9,
    output      wire                        merge_valid_o_7_9,
    input       wire                        merge_ready_i_7_9,
    input       wire        [`DW-1:0]       merge_data_i_7_10,
    input       wire                        merge_valid_i_7_10,
    output      wire                        merge_ready_o_7_10,

    output      wire        [`DW-1:0]       merge_data_o_7_10,
    output      wire                        merge_valid_o_7_10,
    input       wire                        merge_ready_i_7_10,
    input       wire        [`DW-1:0]       merge_data_i_7_11,
    input       wire                        merge_valid_i_7_11,
    output      wire                        merge_ready_o_7_11,

    output      wire        [`DW-1:0]       merge_data_o_7_11,
    output      wire                        merge_valid_o_7_11,
    input       wire                        merge_ready_i_7_11,
    input       wire        [`DW-1:0]       merge_data_i_7_12,
    input       wire                        merge_valid_i_7_12,
    output      wire                        merge_ready_o_7_12,

    output      wire        [`DW-1:0]       merge_data_o_7_12,
    output      wire                        merge_valid_o_7_12,
    input       wire                        merge_ready_i_7_12,
    input       wire        [`DW-1:0]       merge_data_i_7_13,
    input       wire                        merge_valid_i_7_13,
    output      wire                        merge_ready_o_7_13,

    output      wire        [`DW-1:0]       merge_data_o_7_13,
    output      wire                        merge_valid_o_7_13,
    input       wire                        merge_ready_i_7_13,
    input       wire        [`DW-1:0]       merge_data_i_7_14,
    input       wire                        merge_valid_i_7_14,
    output      wire                        merge_ready_o_7_14,

    output      wire        [`DW-1:0]       merge_data_o_7_14,
    output      wire                        merge_valid_o_7_14,
    input       wire                        merge_ready_i_7_14,
    input       wire        [`DW-1:0]       merge_data_i_7_15,
    input       wire                        merge_valid_i_7_15,
    output      wire                        merge_ready_o_7_15,

    output      wire        [`DW-1:0]       merge_data_o_7_15,
    output      wire                        merge_valid_o_7_15,
    input       wire                        merge_ready_i_7_15,
    input       wire        [`DW-1:0]       merge_data_i_7_16,
    input       wire                        merge_valid_i_7_16,
    output      wire                        merge_ready_o_7_16,

    output      wire        [`DW-1:0]       merge_data_o_7_16,
    output      wire                        merge_valid_o_7_16,
    input       wire                        merge_ready_i_7_16,
    input       wire        [`DW-1:0]       merge_data_i_7_17,
    input       wire                        merge_valid_i_7_17,
    output      wire                        merge_ready_o_7_17,

    output      wire        [`DW-1:0]       merge_data_o_7_17,
    output      wire                        merge_valid_o_7_17,
    input       wire                        merge_ready_i_7_17,
    input       wire        [`DW-1:0]       merge_data_i_7_18,
    input       wire                        merge_valid_i_7_18,
    output      wire                        merge_ready_o_7_18,

    output      wire        [`DW-1:0]       merge_data_o_7_18,
    output      wire                        merge_valid_o_7_18,
    input       wire                        merge_ready_i_7_18,
    input       wire        [`DW-1:0]       merge_data_i_7_19,
    input       wire                        merge_valid_i_7_19,
    output      wire                        merge_ready_o_7_19,

    output      wire        [`DW-1:0]       merge_data_o_7_19,
    output      wire                        merge_valid_o_7_19,
    input       wire                        merge_ready_i_7_19,
    input       wire        [`DW-1:0]       merge_data_i_7_20,
    input       wire                        merge_valid_i_7_20,
    output      wire                        merge_ready_o_7_20,

    output      wire        [`DW-1:0]       merge_data_o_7_20,
    output      wire                        merge_valid_o_7_20,
    input       wire                        merge_ready_i_7_20,
    input       wire        [`DW-1:0]       merge_data_i_7_21,
    input       wire                        merge_valid_i_7_21,
    output      wire                        merge_ready_o_7_21,

    output      wire        [`DW-1:0]       merge_data_o_7_21,
    output      wire                        merge_valid_o_7_21,
    input       wire                        merge_ready_i_7_21,
    input       wire        [`DW-1:0]       merge_data_i_7_22,
    input       wire                        merge_valid_i_7_22,
    output      wire                        merge_ready_o_7_22,

    output      wire        [`DW-1:0]       merge_data_o_7_22,
    output      wire                        merge_valid_o_7_22,
    input       wire                        merge_ready_i_7_22,
    input       wire        [`DW-1:0]       merge_data_i_7_23,
    input       wire                        merge_valid_i_7_23,
    output      wire                        merge_ready_o_7_23,

    output      wire        [`DW-1:0]       merge_data_o_7_23,
    output      wire                        merge_valid_o_7_23,
    input       wire                        merge_ready_i_7_23,
    input       wire        [`DW-1:0]       merge_data_i_7_24,
    input       wire                        merge_valid_i_7_24,
    output      wire                        merge_ready_o_7_24,

    output      wire        [`DW-1:0]       merge_data_o_7_24,
    output      wire                        merge_valid_o_7_24,
    input       wire                        merge_ready_i_7_24,
    input       wire        [`DW-1:0]       merge_data_i_8_0,
    input       wire                        merge_valid_i_8_0,
    output      wire                        merge_ready_o_8_0,

    output      wire        [`DW-1:0]       merge_data_o_8_0,
    output      wire                        merge_valid_o_8_0,
    input       wire                        merge_ready_i_8_0,
    input       wire        [`DW-1:0]       merge_data_i_8_1,
    input       wire                        merge_valid_i_8_1,
    output      wire                        merge_ready_o_8_1,

    output      wire        [`DW-1:0]       merge_data_o_8_1,
    output      wire                        merge_valid_o_8_1,
    input       wire                        merge_ready_i_8_1,
    input       wire        [`DW-1:0]       merge_data_i_8_2,
    input       wire                        merge_valid_i_8_2,
    output      wire                        merge_ready_o_8_2,

    output      wire        [`DW-1:0]       merge_data_o_8_2,
    output      wire                        merge_valid_o_8_2,
    input       wire                        merge_ready_i_8_2,
    input       wire        [`DW-1:0]       merge_data_i_8_3,
    input       wire                        merge_valid_i_8_3,
    output      wire                        merge_ready_o_8_3,

    output      wire        [`DW-1:0]       merge_data_o_8_3,
    output      wire                        merge_valid_o_8_3,
    input       wire                        merge_ready_i_8_3,
    input       wire        [`DW-1:0]       merge_data_i_8_4,
    input       wire                        merge_valid_i_8_4,
    output      wire                        merge_ready_o_8_4,

    output      wire        [`DW-1:0]       merge_data_o_8_4,
    output      wire                        merge_valid_o_8_4,
    input       wire                        merge_ready_i_8_4,
    input       wire        [`DW-1:0]       merge_data_i_8_5,
    input       wire                        merge_valid_i_8_5,
    output      wire                        merge_ready_o_8_5,

    output      wire        [`DW-1:0]       merge_data_o_8_5,
    output      wire                        merge_valid_o_8_5,
    input       wire                        merge_ready_i_8_5,
    input       wire        [`DW-1:0]       merge_data_i_8_6,
    input       wire                        merge_valid_i_8_6,
    output      wire                        merge_ready_o_8_6,

    output      wire        [`DW-1:0]       merge_data_o_8_6,
    output      wire                        merge_valid_o_8_6,
    input       wire                        merge_ready_i_8_6,
    input       wire        [`DW-1:0]       merge_data_i_8_7,
    input       wire                        merge_valid_i_8_7,
    output      wire                        merge_ready_o_8_7,

    output      wire        [`DW-1:0]       merge_data_o_8_7,
    output      wire                        merge_valid_o_8_7,
    input       wire                        merge_ready_i_8_7,
    input       wire        [`DW-1:0]       merge_data_i_8_8,
    input       wire                        merge_valid_i_8_8,
    output      wire                        merge_ready_o_8_8,

    output      wire        [`DW-1:0]       merge_data_o_8_8,
    output      wire                        merge_valid_o_8_8,
    input       wire                        merge_ready_i_8_8,
    input       wire        [`DW-1:0]       merge_data_i_8_9,
    input       wire                        merge_valid_i_8_9,
    output      wire                        merge_ready_o_8_9,

    output      wire        [`DW-1:0]       merge_data_o_8_9,
    output      wire                        merge_valid_o_8_9,
    input       wire                        merge_ready_i_8_9,
    input       wire        [`DW-1:0]       merge_data_i_8_10,
    input       wire                        merge_valid_i_8_10,
    output      wire                        merge_ready_o_8_10,

    output      wire        [`DW-1:0]       merge_data_o_8_10,
    output      wire                        merge_valid_o_8_10,
    input       wire                        merge_ready_i_8_10,
    input       wire        [`DW-1:0]       merge_data_i_8_11,
    input       wire                        merge_valid_i_8_11,
    output      wire                        merge_ready_o_8_11,

    output      wire        [`DW-1:0]       merge_data_o_8_11,
    output      wire                        merge_valid_o_8_11,
    input       wire                        merge_ready_i_8_11,
    input       wire        [`DW-1:0]       merge_data_i_8_12,
    input       wire                        merge_valid_i_8_12,
    output      wire                        merge_ready_o_8_12,

    output      wire        [`DW-1:0]       merge_data_o_8_12,
    output      wire                        merge_valid_o_8_12,
    input       wire                        merge_ready_i_8_12,
    input       wire        [`DW-1:0]       merge_data_i_8_13,
    input       wire                        merge_valid_i_8_13,
    output      wire                        merge_ready_o_8_13,

    output      wire        [`DW-1:0]       merge_data_o_8_13,
    output      wire                        merge_valid_o_8_13,
    input       wire                        merge_ready_i_8_13,
    input       wire        [`DW-1:0]       merge_data_i_8_14,
    input       wire                        merge_valid_i_8_14,
    output      wire                        merge_ready_o_8_14,

    output      wire        [`DW-1:0]       merge_data_o_8_14,
    output      wire                        merge_valid_o_8_14,
    input       wire                        merge_ready_i_8_14,
    input       wire        [`DW-1:0]       merge_data_i_8_15,
    input       wire                        merge_valid_i_8_15,
    output      wire                        merge_ready_o_8_15,

    output      wire        [`DW-1:0]       merge_data_o_8_15,
    output      wire                        merge_valid_o_8_15,
    input       wire                        merge_ready_i_8_15,
    input       wire        [`DW-1:0]       merge_data_i_8_16,
    input       wire                        merge_valid_i_8_16,
    output      wire                        merge_ready_o_8_16,

    output      wire        [`DW-1:0]       merge_data_o_8_16,
    output      wire                        merge_valid_o_8_16,
    input       wire                        merge_ready_i_8_16,
    input       wire        [`DW-1:0]       merge_data_i_8_17,
    input       wire                        merge_valid_i_8_17,
    output      wire                        merge_ready_o_8_17,

    output      wire        [`DW-1:0]       merge_data_o_8_17,
    output      wire                        merge_valid_o_8_17,
    input       wire                        merge_ready_i_8_17,
    input       wire        [`DW-1:0]       merge_data_i_8_18,
    input       wire                        merge_valid_i_8_18,
    output      wire                        merge_ready_o_8_18,

    output      wire        [`DW-1:0]       merge_data_o_8_18,
    output      wire                        merge_valid_o_8_18,
    input       wire                        merge_ready_i_8_18,
    input       wire        [`DW-1:0]       merge_data_i_8_19,
    input       wire                        merge_valid_i_8_19,
    output      wire                        merge_ready_o_8_19,

    output      wire        [`DW-1:0]       merge_data_o_8_19,
    output      wire                        merge_valid_o_8_19,
    input       wire                        merge_ready_i_8_19,
    input       wire        [`DW-1:0]       merge_data_i_8_20,
    input       wire                        merge_valid_i_8_20,
    output      wire                        merge_ready_o_8_20,

    output      wire        [`DW-1:0]       merge_data_o_8_20,
    output      wire                        merge_valid_o_8_20,
    input       wire                        merge_ready_i_8_20,
    input       wire        [`DW-1:0]       merge_data_i_8_21,
    input       wire                        merge_valid_i_8_21,
    output      wire                        merge_ready_o_8_21,

    output      wire        [`DW-1:0]       merge_data_o_8_21,
    output      wire                        merge_valid_o_8_21,
    input       wire                        merge_ready_i_8_21,
    input       wire        [`DW-1:0]       merge_data_i_8_22,
    input       wire                        merge_valid_i_8_22,
    output      wire                        merge_ready_o_8_22,

    output      wire        [`DW-1:0]       merge_data_o_8_22,
    output      wire                        merge_valid_o_8_22,
    input       wire                        merge_ready_i_8_22,
    input       wire        [`DW-1:0]       merge_data_i_8_23,
    input       wire                        merge_valid_i_8_23,
    output      wire                        merge_ready_o_8_23,

    output      wire        [`DW-1:0]       merge_data_o_8_23,
    output      wire                        merge_valid_o_8_23,
    input       wire                        merge_ready_i_8_23,
    input       wire        [`DW-1:0]       merge_data_i_8_24,
    input       wire                        merge_valid_i_8_24,
    output      wire                        merge_ready_o_8_24,

    output      wire        [`DW-1:0]       merge_data_o_8_24,
    output      wire                        merge_valid_o_8_24,
    input       wire                        merge_ready_i_8_24,
    input       wire        [`DW-1:0]       merge_data_i_9_0,
    input       wire                        merge_valid_i_9_0,
    output      wire                        merge_ready_o_9_0,

    output      wire        [`DW-1:0]       merge_data_o_9_0,
    output      wire                        merge_valid_o_9_0,
    input       wire                        merge_ready_i_9_0,
    input       wire        [`DW-1:0]       merge_data_i_9_1,
    input       wire                        merge_valid_i_9_1,
    output      wire                        merge_ready_o_9_1,

    output      wire        [`DW-1:0]       merge_data_o_9_1,
    output      wire                        merge_valid_o_9_1,
    input       wire                        merge_ready_i_9_1,
    input       wire        [`DW-1:0]       merge_data_i_9_2,
    input       wire                        merge_valid_i_9_2,
    output      wire                        merge_ready_o_9_2,

    output      wire        [`DW-1:0]       merge_data_o_9_2,
    output      wire                        merge_valid_o_9_2,
    input       wire                        merge_ready_i_9_2,
    input       wire        [`DW-1:0]       merge_data_i_9_3,
    input       wire                        merge_valid_i_9_3,
    output      wire                        merge_ready_o_9_3,

    output      wire        [`DW-1:0]       merge_data_o_9_3,
    output      wire                        merge_valid_o_9_3,
    input       wire                        merge_ready_i_9_3,
    input       wire        [`DW-1:0]       merge_data_i_9_4,
    input       wire                        merge_valid_i_9_4,
    output      wire                        merge_ready_o_9_4,

    output      wire        [`DW-1:0]       merge_data_o_9_4,
    output      wire                        merge_valid_o_9_4,
    input       wire                        merge_ready_i_9_4,
    input       wire        [`DW-1:0]       merge_data_i_9_5,
    input       wire                        merge_valid_i_9_5,
    output      wire                        merge_ready_o_9_5,

    output      wire        [`DW-1:0]       merge_data_o_9_5,
    output      wire                        merge_valid_o_9_5,
    input       wire                        merge_ready_i_9_5,
    input       wire        [`DW-1:0]       merge_data_i_9_6,
    input       wire                        merge_valid_i_9_6,
    output      wire                        merge_ready_o_9_6,

    output      wire        [`DW-1:0]       merge_data_o_9_6,
    output      wire                        merge_valid_o_9_6,
    input       wire                        merge_ready_i_9_6,
    input       wire        [`DW-1:0]       merge_data_i_9_7,
    input       wire                        merge_valid_i_9_7,
    output      wire                        merge_ready_o_9_7,

    output      wire        [`DW-1:0]       merge_data_o_9_7,
    output      wire                        merge_valid_o_9_7,
    input       wire                        merge_ready_i_9_7,
    input       wire        [`DW-1:0]       merge_data_i_9_8,
    input       wire                        merge_valid_i_9_8,
    output      wire                        merge_ready_o_9_8,

    output      wire        [`DW-1:0]       merge_data_o_9_8,
    output      wire                        merge_valid_o_9_8,
    input       wire                        merge_ready_i_9_8,
    input       wire        [`DW-1:0]       merge_data_i_9_9,
    input       wire                        merge_valid_i_9_9,
    output      wire                        merge_ready_o_9_9,

    output      wire        [`DW-1:0]       merge_data_o_9_9,
    output      wire                        merge_valid_o_9_9,
    input       wire                        merge_ready_i_9_9,
    input       wire        [`DW-1:0]       merge_data_i_9_10,
    input       wire                        merge_valid_i_9_10,
    output      wire                        merge_ready_o_9_10,

    output      wire        [`DW-1:0]       merge_data_o_9_10,
    output      wire                        merge_valid_o_9_10,
    input       wire                        merge_ready_i_9_10,
    input       wire        [`DW-1:0]       merge_data_i_9_11,
    input       wire                        merge_valid_i_9_11,
    output      wire                        merge_ready_o_9_11,

    output      wire        [`DW-1:0]       merge_data_o_9_11,
    output      wire                        merge_valid_o_9_11,
    input       wire                        merge_ready_i_9_11,
    input       wire        [`DW-1:0]       merge_data_i_9_12,
    input       wire                        merge_valid_i_9_12,
    output      wire                        merge_ready_o_9_12,

    output      wire        [`DW-1:0]       merge_data_o_9_12,
    output      wire                        merge_valid_o_9_12,
    input       wire                        merge_ready_i_9_12,
    input       wire        [`DW-1:0]       merge_data_i_9_13,
    input       wire                        merge_valid_i_9_13,
    output      wire                        merge_ready_o_9_13,

    output      wire        [`DW-1:0]       merge_data_o_9_13,
    output      wire                        merge_valid_o_9_13,
    input       wire                        merge_ready_i_9_13,
    input       wire        [`DW-1:0]       merge_data_i_9_14,
    input       wire                        merge_valid_i_9_14,
    output      wire                        merge_ready_o_9_14,

    output      wire        [`DW-1:0]       merge_data_o_9_14,
    output      wire                        merge_valid_o_9_14,
    input       wire                        merge_ready_i_9_14,
    input       wire        [`DW-1:0]       merge_data_i_9_15,
    input       wire                        merge_valid_i_9_15,
    output      wire                        merge_ready_o_9_15,

    output      wire        [`DW-1:0]       merge_data_o_9_15,
    output      wire                        merge_valid_o_9_15,
    input       wire                        merge_ready_i_9_15,
    input       wire        [`DW-1:0]       merge_data_i_9_16,
    input       wire                        merge_valid_i_9_16,
    output      wire                        merge_ready_o_9_16,

    output      wire        [`DW-1:0]       merge_data_o_9_16,
    output      wire                        merge_valid_o_9_16,
    input       wire                        merge_ready_i_9_16,
    input       wire        [`DW-1:0]       merge_data_i_9_17,
    input       wire                        merge_valid_i_9_17,
    output      wire                        merge_ready_o_9_17,

    output      wire        [`DW-1:0]       merge_data_o_9_17,
    output      wire                        merge_valid_o_9_17,
    input       wire                        merge_ready_i_9_17,
    input       wire        [`DW-1:0]       merge_data_i_9_18,
    input       wire                        merge_valid_i_9_18,
    output      wire                        merge_ready_o_9_18,

    output      wire        [`DW-1:0]       merge_data_o_9_18,
    output      wire                        merge_valid_o_9_18,
    input       wire                        merge_ready_i_9_18,
    input       wire        [`DW-1:0]       merge_data_i_9_19,
    input       wire                        merge_valid_i_9_19,
    output      wire                        merge_ready_o_9_19,

    output      wire        [`DW-1:0]       merge_data_o_9_19,
    output      wire                        merge_valid_o_9_19,
    input       wire                        merge_ready_i_9_19,
    input       wire        [`DW-1:0]       merge_data_i_9_20,
    input       wire                        merge_valid_i_9_20,
    output      wire                        merge_ready_o_9_20,

    output      wire        [`DW-1:0]       merge_data_o_9_20,
    output      wire                        merge_valid_o_9_20,
    input       wire                        merge_ready_i_9_20,
    input       wire        [`DW-1:0]       merge_data_i_9_21,
    input       wire                        merge_valid_i_9_21,
    output      wire                        merge_ready_o_9_21,

    output      wire        [`DW-1:0]       merge_data_o_9_21,
    output      wire                        merge_valid_o_9_21,
    input       wire                        merge_ready_i_9_21,
    input       wire        [`DW-1:0]       merge_data_i_9_22,
    input       wire                        merge_valid_i_9_22,
    output      wire                        merge_ready_o_9_22,

    output      wire        [`DW-1:0]       merge_data_o_9_22,
    output      wire                        merge_valid_o_9_22,
    input       wire                        merge_ready_i_9_22,
    input       wire        [`DW-1:0]       merge_data_i_9_23,
    input       wire                        merge_valid_i_9_23,
    output      wire                        merge_ready_o_9_23,

    output      wire        [`DW-1:0]       merge_data_o_9_23,
    output      wire                        merge_valid_o_9_23,
    input       wire                        merge_ready_i_9_23,
    input       wire        [`DW-1:0]       merge_data_i_9_24,
    input       wire                        merge_valid_i_9_24,
    output      wire                        merge_ready_o_9_24,

    output      wire        [`DW-1:0]       merge_data_o_9_24,
    output      wire                        merge_valid_o_9_24,
    input       wire                        merge_ready_i_9_24,
    input       wire        [`DW-1:0]       gather_data_i_0_0,
    input       wire                        gather_valid_i_0_0,
    output      wire                        gather_ready_o_0_0,

    output      wire        [`DW-1:0]       gather_data_o_0_0,
    output      wire                        gather_valid_o_0_0,
    input       wire                        gather_ready_i_0_0,
    input       wire        [`DW-1:0]       gather_data_i_0_1,
    input       wire                        gather_valid_i_0_1,
    output      wire                        gather_ready_o_0_1,

    output      wire        [`DW-1:0]       gather_data_o_0_1,
    output      wire                        gather_valid_o_0_1,
    input       wire                        gather_ready_i_0_1,
    input       wire        [`DW-1:0]       gather_data_i_0_2,
    input       wire                        gather_valid_i_0_2,
    output      wire                        gather_ready_o_0_2,

    output      wire        [`DW-1:0]       gather_data_o_0_2,
    output      wire                        gather_valid_o_0_2,
    input       wire                        gather_ready_i_0_2,
    input       wire        [`DW-1:0]       gather_data_i_0_3,
    input       wire                        gather_valid_i_0_3,
    output      wire                        gather_ready_o_0_3,

    output      wire        [`DW-1:0]       gather_data_o_0_3,
    output      wire                        gather_valid_o_0_3,
    input       wire                        gather_ready_i_0_3,
    input       wire        [`DW-1:0]       gather_data_i_0_4,
    input       wire                        gather_valid_i_0_4,
    output      wire                        gather_ready_o_0_4,

    output      wire        [`DW-1:0]       gather_data_o_0_4,
    output      wire                        gather_valid_o_0_4,
    input       wire                        gather_ready_i_0_4,
    input       wire        [`DW-1:0]       gather_data_i_0_5,
    input       wire                        gather_valid_i_0_5,
    output      wire                        gather_ready_o_0_5,

    output      wire        [`DW-1:0]       gather_data_o_0_5,
    output      wire                        gather_valid_o_0_5,
    input       wire                        gather_ready_i_0_5,
    input       wire        [`DW-1:0]       gather_data_i_0_6,
    input       wire                        gather_valid_i_0_6,
    output      wire                        gather_ready_o_0_6,

    output      wire        [`DW-1:0]       gather_data_o_0_6,
    output      wire                        gather_valid_o_0_6,
    input       wire                        gather_ready_i_0_6,
    input       wire        [`DW-1:0]       gather_data_i_0_7,
    input       wire                        gather_valid_i_0_7,
    output      wire                        gather_ready_o_0_7,

    output      wire        [`DW-1:0]       gather_data_o_0_7,
    output      wire                        gather_valid_o_0_7,
    input       wire                        gather_ready_i_0_7,
    input       wire        [`DW-1:0]       gather_data_i_0_8,
    input       wire                        gather_valid_i_0_8,
    output      wire                        gather_ready_o_0_8,

    output      wire        [`DW-1:0]       gather_data_o_0_8,
    output      wire                        gather_valid_o_0_8,
    input       wire                        gather_ready_i_0_8,
    input       wire        [`DW-1:0]       gather_data_i_0_9,
    input       wire                        gather_valid_i_0_9,
    output      wire                        gather_ready_o_0_9,

    output      wire        [`DW-1:0]       gather_data_o_0_9,
    output      wire                        gather_valid_o_0_9,
    input       wire                        gather_ready_i_0_9,
    input       wire        [`DW-1:0]       gather_data_i_0_10,
    input       wire                        gather_valid_i_0_10,
    output      wire                        gather_ready_o_0_10,

    output      wire        [`DW-1:0]       gather_data_o_0_10,
    output      wire                        gather_valid_o_0_10,
    input       wire                        gather_ready_i_0_10,
    input       wire        [`DW-1:0]       gather_data_i_0_11,
    input       wire                        gather_valid_i_0_11,
    output      wire                        gather_ready_o_0_11,

    output      wire        [`DW-1:0]       gather_data_o_0_11,
    output      wire                        gather_valid_o_0_11,
    input       wire                        gather_ready_i_0_11,
    input       wire        [`DW-1:0]       gather_data_i_0_12,
    input       wire                        gather_valid_i_0_12,
    output      wire                        gather_ready_o_0_12,

    output      wire        [`DW-1:0]       gather_data_o_0_12,
    output      wire                        gather_valid_o_0_12,
    input       wire                        gather_ready_i_0_12,
    input       wire        [`DW-1:0]       gather_data_i_0_13,
    input       wire                        gather_valid_i_0_13,
    output      wire                        gather_ready_o_0_13,

    output      wire        [`DW-1:0]       gather_data_o_0_13,
    output      wire                        gather_valid_o_0_13,
    input       wire                        gather_ready_i_0_13,
    input       wire        [`DW-1:0]       gather_data_i_0_14,
    input       wire                        gather_valid_i_0_14,
    output      wire                        gather_ready_o_0_14,

    output      wire        [`DW-1:0]       gather_data_o_0_14,
    output      wire                        gather_valid_o_0_14,
    input       wire                        gather_ready_i_0_14,
    input       wire        [`DW-1:0]       gather_data_i_0_15,
    input       wire                        gather_valid_i_0_15,
    output      wire                        gather_ready_o_0_15,

    output      wire        [`DW-1:0]       gather_data_o_0_15,
    output      wire                        gather_valid_o_0_15,
    input       wire                        gather_ready_i_0_15,
    input       wire        [`DW-1:0]       gather_data_i_0_16,
    input       wire                        gather_valid_i_0_16,
    output      wire                        gather_ready_o_0_16,

    output      wire        [`DW-1:0]       gather_data_o_0_16,
    output      wire                        gather_valid_o_0_16,
    input       wire                        gather_ready_i_0_16,
    input       wire        [`DW-1:0]       gather_data_i_0_17,
    input       wire                        gather_valid_i_0_17,
    output      wire                        gather_ready_o_0_17,

    output      wire        [`DW-1:0]       gather_data_o_0_17,
    output      wire                        gather_valid_o_0_17,
    input       wire                        gather_ready_i_0_17,
    input       wire        [`DW-1:0]       gather_data_i_0_18,
    input       wire                        gather_valid_i_0_18,
    output      wire                        gather_ready_o_0_18,

    output      wire        [`DW-1:0]       gather_data_o_0_18,
    output      wire                        gather_valid_o_0_18,
    input       wire                        gather_ready_i_0_18,
    input       wire        [`DW-1:0]       gather_data_i_0_19,
    input       wire                        gather_valid_i_0_19,
    output      wire                        gather_ready_o_0_19,

    output      wire        [`DW-1:0]       gather_data_o_0_19,
    output      wire                        gather_valid_o_0_19,
    input       wire                        gather_ready_i_0_19,
    input       wire        [`DW-1:0]       gather_data_i_0_20,
    input       wire                        gather_valid_i_0_20,
    output      wire                        gather_ready_o_0_20,

    output      wire        [`DW-1:0]       gather_data_o_0_20,
    output      wire                        gather_valid_o_0_20,
    input       wire                        gather_ready_i_0_20,
    input       wire        [`DW-1:0]       gather_data_i_0_21,
    input       wire                        gather_valid_i_0_21,
    output      wire                        gather_ready_o_0_21,

    output      wire        [`DW-1:0]       gather_data_o_0_21,
    output      wire                        gather_valid_o_0_21,
    input       wire                        gather_ready_i_0_21,
    input       wire        [`DW-1:0]       gather_data_i_0_22,
    input       wire                        gather_valid_i_0_22,
    output      wire                        gather_ready_o_0_22,

    output      wire        [`DW-1:0]       gather_data_o_0_22,
    output      wire                        gather_valid_o_0_22,
    input       wire                        gather_ready_i_0_22,
    input       wire        [`DW-1:0]       gather_data_i_0_23,
    input       wire                        gather_valid_i_0_23,
    output      wire                        gather_ready_o_0_23,

    output      wire        [`DW-1:0]       gather_data_o_0_23,
    output      wire                        gather_valid_o_0_23,
    input       wire                        gather_ready_i_0_23,
    input       wire        [`DW-1:0]       gather_data_i_0_24,
    input       wire                        gather_valid_i_0_24,
    output      wire                        gather_ready_o_0_24,

    output      wire        [`DW-1:0]       gather_data_o_0_24,
    output      wire                        gather_valid_o_0_24,
    input       wire                        gather_ready_i_0_24,
    input       wire        [`DW-1:0]       gather_data_i_1_0,
    input       wire                        gather_valid_i_1_0,
    output      wire                        gather_ready_o_1_0,

    output      wire        [`DW-1:0]       gather_data_o_1_0,
    output      wire                        gather_valid_o_1_0,
    input       wire                        gather_ready_i_1_0,
    input       wire        [`DW-1:0]       gather_data_i_1_1,
    input       wire                        gather_valid_i_1_1,
    output      wire                        gather_ready_o_1_1,

    output      wire        [`DW-1:0]       gather_data_o_1_1,
    output      wire                        gather_valid_o_1_1,
    input       wire                        gather_ready_i_1_1,
    input       wire        [`DW-1:0]       gather_data_i_1_2,
    input       wire                        gather_valid_i_1_2,
    output      wire                        gather_ready_o_1_2,

    output      wire        [`DW-1:0]       gather_data_o_1_2,
    output      wire                        gather_valid_o_1_2,
    input       wire                        gather_ready_i_1_2,
    input       wire        [`DW-1:0]       gather_data_i_1_3,
    input       wire                        gather_valid_i_1_3,
    output      wire                        gather_ready_o_1_3,

    output      wire        [`DW-1:0]       gather_data_o_1_3,
    output      wire                        gather_valid_o_1_3,
    input       wire                        gather_ready_i_1_3,
    input       wire        [`DW-1:0]       gather_data_i_1_4,
    input       wire                        gather_valid_i_1_4,
    output      wire                        gather_ready_o_1_4,

    output      wire        [`DW-1:0]       gather_data_o_1_4,
    output      wire                        gather_valid_o_1_4,
    input       wire                        gather_ready_i_1_4,
    input       wire        [`DW-1:0]       gather_data_i_1_5,
    input       wire                        gather_valid_i_1_5,
    output      wire                        gather_ready_o_1_5,

    output      wire        [`DW-1:0]       gather_data_o_1_5,
    output      wire                        gather_valid_o_1_5,
    input       wire                        gather_ready_i_1_5,
    input       wire        [`DW-1:0]       gather_data_i_1_6,
    input       wire                        gather_valid_i_1_6,
    output      wire                        gather_ready_o_1_6,

    output      wire        [`DW-1:0]       gather_data_o_1_6,
    output      wire                        gather_valid_o_1_6,
    input       wire                        gather_ready_i_1_6,
    input       wire        [`DW-1:0]       gather_data_i_1_7,
    input       wire                        gather_valid_i_1_7,
    output      wire                        gather_ready_o_1_7,

    output      wire        [`DW-1:0]       gather_data_o_1_7,
    output      wire                        gather_valid_o_1_7,
    input       wire                        gather_ready_i_1_7,
    input       wire        [`DW-1:0]       gather_data_i_1_8,
    input       wire                        gather_valid_i_1_8,
    output      wire                        gather_ready_o_1_8,

    output      wire        [`DW-1:0]       gather_data_o_1_8,
    output      wire                        gather_valid_o_1_8,
    input       wire                        gather_ready_i_1_8,
    input       wire        [`DW-1:0]       gather_data_i_1_9,
    input       wire                        gather_valid_i_1_9,
    output      wire                        gather_ready_o_1_9,

    output      wire        [`DW-1:0]       gather_data_o_1_9,
    output      wire                        gather_valid_o_1_9,
    input       wire                        gather_ready_i_1_9,
    input       wire        [`DW-1:0]       gather_data_i_1_10,
    input       wire                        gather_valid_i_1_10,
    output      wire                        gather_ready_o_1_10,

    output      wire        [`DW-1:0]       gather_data_o_1_10,
    output      wire                        gather_valid_o_1_10,
    input       wire                        gather_ready_i_1_10,
    input       wire        [`DW-1:0]       gather_data_i_1_11,
    input       wire                        gather_valid_i_1_11,
    output      wire                        gather_ready_o_1_11,

    output      wire        [`DW-1:0]       gather_data_o_1_11,
    output      wire                        gather_valid_o_1_11,
    input       wire                        gather_ready_i_1_11,
    input       wire        [`DW-1:0]       gather_data_i_1_12,
    input       wire                        gather_valid_i_1_12,
    output      wire                        gather_ready_o_1_12,

    output      wire        [`DW-1:0]       gather_data_o_1_12,
    output      wire                        gather_valid_o_1_12,
    input       wire                        gather_ready_i_1_12,
    input       wire        [`DW-1:0]       gather_data_i_1_13,
    input       wire                        gather_valid_i_1_13,
    output      wire                        gather_ready_o_1_13,

    output      wire        [`DW-1:0]       gather_data_o_1_13,
    output      wire                        gather_valid_o_1_13,
    input       wire                        gather_ready_i_1_13,
    input       wire        [`DW-1:0]       gather_data_i_1_14,
    input       wire                        gather_valid_i_1_14,
    output      wire                        gather_ready_o_1_14,

    output      wire        [`DW-1:0]       gather_data_o_1_14,
    output      wire                        gather_valid_o_1_14,
    input       wire                        gather_ready_i_1_14,
    input       wire        [`DW-1:0]       gather_data_i_1_15,
    input       wire                        gather_valid_i_1_15,
    output      wire                        gather_ready_o_1_15,

    output      wire        [`DW-1:0]       gather_data_o_1_15,
    output      wire                        gather_valid_o_1_15,
    input       wire                        gather_ready_i_1_15,
    input       wire        [`DW-1:0]       gather_data_i_1_16,
    input       wire                        gather_valid_i_1_16,
    output      wire                        gather_ready_o_1_16,

    output      wire        [`DW-1:0]       gather_data_o_1_16,
    output      wire                        gather_valid_o_1_16,
    input       wire                        gather_ready_i_1_16,
    input       wire        [`DW-1:0]       gather_data_i_1_17,
    input       wire                        gather_valid_i_1_17,
    output      wire                        gather_ready_o_1_17,

    output      wire        [`DW-1:0]       gather_data_o_1_17,
    output      wire                        gather_valid_o_1_17,
    input       wire                        gather_ready_i_1_17,
    input       wire        [`DW-1:0]       gather_data_i_1_18,
    input       wire                        gather_valid_i_1_18,
    output      wire                        gather_ready_o_1_18,

    output      wire        [`DW-1:0]       gather_data_o_1_18,
    output      wire                        gather_valid_o_1_18,
    input       wire                        gather_ready_i_1_18,
    input       wire        [`DW-1:0]       gather_data_i_1_19,
    input       wire                        gather_valid_i_1_19,
    output      wire                        gather_ready_o_1_19,

    output      wire        [`DW-1:0]       gather_data_o_1_19,
    output      wire                        gather_valid_o_1_19,
    input       wire                        gather_ready_i_1_19,
    input       wire        [`DW-1:0]       gather_data_i_1_20,
    input       wire                        gather_valid_i_1_20,
    output      wire                        gather_ready_o_1_20,

    output      wire        [`DW-1:0]       gather_data_o_1_20,
    output      wire                        gather_valid_o_1_20,
    input       wire                        gather_ready_i_1_20,
    input       wire        [`DW-1:0]       gather_data_i_1_21,
    input       wire                        gather_valid_i_1_21,
    output      wire                        gather_ready_o_1_21,

    output      wire        [`DW-1:0]       gather_data_o_1_21,
    output      wire                        gather_valid_o_1_21,
    input       wire                        gather_ready_i_1_21,
    input       wire        [`DW-1:0]       gather_data_i_1_22,
    input       wire                        gather_valid_i_1_22,
    output      wire                        gather_ready_o_1_22,

    output      wire        [`DW-1:0]       gather_data_o_1_22,
    output      wire                        gather_valid_o_1_22,
    input       wire                        gather_ready_i_1_22,
    input       wire        [`DW-1:0]       gather_data_i_1_23,
    input       wire                        gather_valid_i_1_23,
    output      wire                        gather_ready_o_1_23,

    output      wire        [`DW-1:0]       gather_data_o_1_23,
    output      wire                        gather_valid_o_1_23,
    input       wire                        gather_ready_i_1_23,
    input       wire        [`DW-1:0]       gather_data_i_1_24,
    input       wire                        gather_valid_i_1_24,
    output      wire                        gather_ready_o_1_24,

    output      wire        [`DW-1:0]       gather_data_o_1_24,
    output      wire                        gather_valid_o_1_24,
    input       wire                        gather_ready_i_1_24,
    input       wire        [`DW-1:0]       gather_data_i_2_0,
    input       wire                        gather_valid_i_2_0,
    output      wire                        gather_ready_o_2_0,

    output      wire        [`DW-1:0]       gather_data_o_2_0,
    output      wire                        gather_valid_o_2_0,
    input       wire                        gather_ready_i_2_0,
    input       wire        [`DW-1:0]       gather_data_i_2_1,
    input       wire                        gather_valid_i_2_1,
    output      wire                        gather_ready_o_2_1,

    output      wire        [`DW-1:0]       gather_data_o_2_1,
    output      wire                        gather_valid_o_2_1,
    input       wire                        gather_ready_i_2_1,
    input       wire        [`DW-1:0]       gather_data_i_2_2,
    input       wire                        gather_valid_i_2_2,
    output      wire                        gather_ready_o_2_2,

    output      wire        [`DW-1:0]       gather_data_o_2_2,
    output      wire                        gather_valid_o_2_2,
    input       wire                        gather_ready_i_2_2,
    input       wire        [`DW-1:0]       gather_data_i_2_3,
    input       wire                        gather_valid_i_2_3,
    output      wire                        gather_ready_o_2_3,

    output      wire        [`DW-1:0]       gather_data_o_2_3,
    output      wire                        gather_valid_o_2_3,
    input       wire                        gather_ready_i_2_3,
    input       wire        [`DW-1:0]       gather_data_i_2_4,
    input       wire                        gather_valid_i_2_4,
    output      wire                        gather_ready_o_2_4,

    output      wire        [`DW-1:0]       gather_data_o_2_4,
    output      wire                        gather_valid_o_2_4,
    input       wire                        gather_ready_i_2_4,
    input       wire        [`DW-1:0]       gather_data_i_2_5,
    input       wire                        gather_valid_i_2_5,
    output      wire                        gather_ready_o_2_5,

    output      wire        [`DW-1:0]       gather_data_o_2_5,
    output      wire                        gather_valid_o_2_5,
    input       wire                        gather_ready_i_2_5,
    input       wire        [`DW-1:0]       gather_data_i_2_6,
    input       wire                        gather_valid_i_2_6,
    output      wire                        gather_ready_o_2_6,

    output      wire        [`DW-1:0]       gather_data_o_2_6,
    output      wire                        gather_valid_o_2_6,
    input       wire                        gather_ready_i_2_6,
    input       wire        [`DW-1:0]       gather_data_i_2_7,
    input       wire                        gather_valid_i_2_7,
    output      wire                        gather_ready_o_2_7,

    output      wire        [`DW-1:0]       gather_data_o_2_7,
    output      wire                        gather_valid_o_2_7,
    input       wire                        gather_ready_i_2_7,
    input       wire        [`DW-1:0]       gather_data_i_2_8,
    input       wire                        gather_valid_i_2_8,
    output      wire                        gather_ready_o_2_8,

    output      wire        [`DW-1:0]       gather_data_o_2_8,
    output      wire                        gather_valid_o_2_8,
    input       wire                        gather_ready_i_2_8,
    input       wire        [`DW-1:0]       gather_data_i_2_9,
    input       wire                        gather_valid_i_2_9,
    output      wire                        gather_ready_o_2_9,

    output      wire        [`DW-1:0]       gather_data_o_2_9,
    output      wire                        gather_valid_o_2_9,
    input       wire                        gather_ready_i_2_9,
    input       wire        [`DW-1:0]       gather_data_i_2_10,
    input       wire                        gather_valid_i_2_10,
    output      wire                        gather_ready_o_2_10,

    output      wire        [`DW-1:0]       gather_data_o_2_10,
    output      wire                        gather_valid_o_2_10,
    input       wire                        gather_ready_i_2_10,
    input       wire        [`DW-1:0]       gather_data_i_2_11,
    input       wire                        gather_valid_i_2_11,
    output      wire                        gather_ready_o_2_11,

    output      wire        [`DW-1:0]       gather_data_o_2_11,
    output      wire                        gather_valid_o_2_11,
    input       wire                        gather_ready_i_2_11,
    input       wire        [`DW-1:0]       gather_data_i_2_12,
    input       wire                        gather_valid_i_2_12,
    output      wire                        gather_ready_o_2_12,

    output      wire        [`DW-1:0]       gather_data_o_2_12,
    output      wire                        gather_valid_o_2_12,
    input       wire                        gather_ready_i_2_12,
    input       wire        [`DW-1:0]       gather_data_i_2_13,
    input       wire                        gather_valid_i_2_13,
    output      wire                        gather_ready_o_2_13,

    output      wire        [`DW-1:0]       gather_data_o_2_13,
    output      wire                        gather_valid_o_2_13,
    input       wire                        gather_ready_i_2_13,
    input       wire        [`DW-1:0]       gather_data_i_2_14,
    input       wire                        gather_valid_i_2_14,
    output      wire                        gather_ready_o_2_14,

    output      wire        [`DW-1:0]       gather_data_o_2_14,
    output      wire                        gather_valid_o_2_14,
    input       wire                        gather_ready_i_2_14,
    input       wire        [`DW-1:0]       gather_data_i_2_15,
    input       wire                        gather_valid_i_2_15,
    output      wire                        gather_ready_o_2_15,

    output      wire        [`DW-1:0]       gather_data_o_2_15,
    output      wire                        gather_valid_o_2_15,
    input       wire                        gather_ready_i_2_15,
    input       wire        [`DW-1:0]       gather_data_i_2_16,
    input       wire                        gather_valid_i_2_16,
    output      wire                        gather_ready_o_2_16,

    output      wire        [`DW-1:0]       gather_data_o_2_16,
    output      wire                        gather_valid_o_2_16,
    input       wire                        gather_ready_i_2_16,
    input       wire        [`DW-1:0]       gather_data_i_2_17,
    input       wire                        gather_valid_i_2_17,
    output      wire                        gather_ready_o_2_17,

    output      wire        [`DW-1:0]       gather_data_o_2_17,
    output      wire                        gather_valid_o_2_17,
    input       wire                        gather_ready_i_2_17,
    input       wire        [`DW-1:0]       gather_data_i_2_18,
    input       wire                        gather_valid_i_2_18,
    output      wire                        gather_ready_o_2_18,

    output      wire        [`DW-1:0]       gather_data_o_2_18,
    output      wire                        gather_valid_o_2_18,
    input       wire                        gather_ready_i_2_18,
    input       wire        [`DW-1:0]       gather_data_i_2_19,
    input       wire                        gather_valid_i_2_19,
    output      wire                        gather_ready_o_2_19,

    output      wire        [`DW-1:0]       gather_data_o_2_19,
    output      wire                        gather_valid_o_2_19,
    input       wire                        gather_ready_i_2_19,
    input       wire        [`DW-1:0]       gather_data_i_2_20,
    input       wire                        gather_valid_i_2_20,
    output      wire                        gather_ready_o_2_20,

    output      wire        [`DW-1:0]       gather_data_o_2_20,
    output      wire                        gather_valid_o_2_20,
    input       wire                        gather_ready_i_2_20,
    input       wire        [`DW-1:0]       gather_data_i_2_21,
    input       wire                        gather_valid_i_2_21,
    output      wire                        gather_ready_o_2_21,

    output      wire        [`DW-1:0]       gather_data_o_2_21,
    output      wire                        gather_valid_o_2_21,
    input       wire                        gather_ready_i_2_21,
    input       wire        [`DW-1:0]       gather_data_i_2_22,
    input       wire                        gather_valid_i_2_22,
    output      wire                        gather_ready_o_2_22,

    output      wire        [`DW-1:0]       gather_data_o_2_22,
    output      wire                        gather_valid_o_2_22,
    input       wire                        gather_ready_i_2_22,
    input       wire        [`DW-1:0]       gather_data_i_2_23,
    input       wire                        gather_valid_i_2_23,
    output      wire                        gather_ready_o_2_23,

    output      wire        [`DW-1:0]       gather_data_o_2_23,
    output      wire                        gather_valid_o_2_23,
    input       wire                        gather_ready_i_2_23,
    input       wire        [`DW-1:0]       gather_data_i_2_24,
    input       wire                        gather_valid_i_2_24,
    output      wire                        gather_ready_o_2_24,

    output      wire        [`DW-1:0]       gather_data_o_2_24,
    output      wire                        gather_valid_o_2_24,
    input       wire                        gather_ready_i_2_24,
    input       wire        [`DW-1:0]       gather_data_i_3_0,
    input       wire                        gather_valid_i_3_0,
    output      wire                        gather_ready_o_3_0,

    output      wire        [`DW-1:0]       gather_data_o_3_0,
    output      wire                        gather_valid_o_3_0,
    input       wire                        gather_ready_i_3_0,
    input       wire        [`DW-1:0]       gather_data_i_3_1,
    input       wire                        gather_valid_i_3_1,
    output      wire                        gather_ready_o_3_1,

    output      wire        [`DW-1:0]       gather_data_o_3_1,
    output      wire                        gather_valid_o_3_1,
    input       wire                        gather_ready_i_3_1,
    input       wire        [`DW-1:0]       gather_data_i_3_2,
    input       wire                        gather_valid_i_3_2,
    output      wire                        gather_ready_o_3_2,

    output      wire        [`DW-1:0]       gather_data_o_3_2,
    output      wire                        gather_valid_o_3_2,
    input       wire                        gather_ready_i_3_2,
    input       wire        [`DW-1:0]       gather_data_i_3_3,
    input       wire                        gather_valid_i_3_3,
    output      wire                        gather_ready_o_3_3,

    output      wire        [`DW-1:0]       gather_data_o_3_3,
    output      wire                        gather_valid_o_3_3,
    input       wire                        gather_ready_i_3_3,
    input       wire        [`DW-1:0]       gather_data_i_3_4,
    input       wire                        gather_valid_i_3_4,
    output      wire                        gather_ready_o_3_4,

    output      wire        [`DW-1:0]       gather_data_o_3_4,
    output      wire                        gather_valid_o_3_4,
    input       wire                        gather_ready_i_3_4,
    input       wire        [`DW-1:0]       gather_data_i_3_5,
    input       wire                        gather_valid_i_3_5,
    output      wire                        gather_ready_o_3_5,

    output      wire        [`DW-1:0]       gather_data_o_3_5,
    output      wire                        gather_valid_o_3_5,
    input       wire                        gather_ready_i_3_5,
    input       wire        [`DW-1:0]       gather_data_i_3_6,
    input       wire                        gather_valid_i_3_6,
    output      wire                        gather_ready_o_3_6,

    output      wire        [`DW-1:0]       gather_data_o_3_6,
    output      wire                        gather_valid_o_3_6,
    input       wire                        gather_ready_i_3_6,
    input       wire        [`DW-1:0]       gather_data_i_3_7,
    input       wire                        gather_valid_i_3_7,
    output      wire                        gather_ready_o_3_7,

    output      wire        [`DW-1:0]       gather_data_o_3_7,
    output      wire                        gather_valid_o_3_7,
    input       wire                        gather_ready_i_3_7,
    input       wire        [`DW-1:0]       gather_data_i_3_8,
    input       wire                        gather_valid_i_3_8,
    output      wire                        gather_ready_o_3_8,

    output      wire        [`DW-1:0]       gather_data_o_3_8,
    output      wire                        gather_valid_o_3_8,
    input       wire                        gather_ready_i_3_8,
    input       wire        [`DW-1:0]       gather_data_i_3_9,
    input       wire                        gather_valid_i_3_9,
    output      wire                        gather_ready_o_3_9,

    output      wire        [`DW-1:0]       gather_data_o_3_9,
    output      wire                        gather_valid_o_3_9,
    input       wire                        gather_ready_i_3_9,
    input       wire        [`DW-1:0]       gather_data_i_3_10,
    input       wire                        gather_valid_i_3_10,
    output      wire                        gather_ready_o_3_10,

    output      wire        [`DW-1:0]       gather_data_o_3_10,
    output      wire                        gather_valid_o_3_10,
    input       wire                        gather_ready_i_3_10,
    input       wire        [`DW-1:0]       gather_data_i_3_11,
    input       wire                        gather_valid_i_3_11,
    output      wire                        gather_ready_o_3_11,

    output      wire        [`DW-1:0]       gather_data_o_3_11,
    output      wire                        gather_valid_o_3_11,
    input       wire                        gather_ready_i_3_11,
    input       wire        [`DW-1:0]       gather_data_i_3_12,
    input       wire                        gather_valid_i_3_12,
    output      wire                        gather_ready_o_3_12,

    output      wire        [`DW-1:0]       gather_data_o_3_12,
    output      wire                        gather_valid_o_3_12,
    input       wire                        gather_ready_i_3_12,
    input       wire        [`DW-1:0]       gather_data_i_3_13,
    input       wire                        gather_valid_i_3_13,
    output      wire                        gather_ready_o_3_13,

    output      wire        [`DW-1:0]       gather_data_o_3_13,
    output      wire                        gather_valid_o_3_13,
    input       wire                        gather_ready_i_3_13,
    input       wire        [`DW-1:0]       gather_data_i_3_14,
    input       wire                        gather_valid_i_3_14,
    output      wire                        gather_ready_o_3_14,

    output      wire        [`DW-1:0]       gather_data_o_3_14,
    output      wire                        gather_valid_o_3_14,
    input       wire                        gather_ready_i_3_14,
    input       wire        [`DW-1:0]       gather_data_i_3_15,
    input       wire                        gather_valid_i_3_15,
    output      wire                        gather_ready_o_3_15,

    output      wire        [`DW-1:0]       gather_data_o_3_15,
    output      wire                        gather_valid_o_3_15,
    input       wire                        gather_ready_i_3_15,
    input       wire        [`DW-1:0]       gather_data_i_3_16,
    input       wire                        gather_valid_i_3_16,
    output      wire                        gather_ready_o_3_16,

    output      wire        [`DW-1:0]       gather_data_o_3_16,
    output      wire                        gather_valid_o_3_16,
    input       wire                        gather_ready_i_3_16,
    input       wire        [`DW-1:0]       gather_data_i_3_17,
    input       wire                        gather_valid_i_3_17,
    output      wire                        gather_ready_o_3_17,

    output      wire        [`DW-1:0]       gather_data_o_3_17,
    output      wire                        gather_valid_o_3_17,
    input       wire                        gather_ready_i_3_17,
    input       wire        [`DW-1:0]       gather_data_i_3_18,
    input       wire                        gather_valid_i_3_18,
    output      wire                        gather_ready_o_3_18,

    output      wire        [`DW-1:0]       gather_data_o_3_18,
    output      wire                        gather_valid_o_3_18,
    input       wire                        gather_ready_i_3_18,
    input       wire        [`DW-1:0]       gather_data_i_3_19,
    input       wire                        gather_valid_i_3_19,
    output      wire                        gather_ready_o_3_19,

    output      wire        [`DW-1:0]       gather_data_o_3_19,
    output      wire                        gather_valid_o_3_19,
    input       wire                        gather_ready_i_3_19,
    input       wire        [`DW-1:0]       gather_data_i_3_20,
    input       wire                        gather_valid_i_3_20,
    output      wire                        gather_ready_o_3_20,

    output      wire        [`DW-1:0]       gather_data_o_3_20,
    output      wire                        gather_valid_o_3_20,
    input       wire                        gather_ready_i_3_20,
    input       wire        [`DW-1:0]       gather_data_i_3_21,
    input       wire                        gather_valid_i_3_21,
    output      wire                        gather_ready_o_3_21,

    output      wire        [`DW-1:0]       gather_data_o_3_21,
    output      wire                        gather_valid_o_3_21,
    input       wire                        gather_ready_i_3_21,
    input       wire        [`DW-1:0]       gather_data_i_3_22,
    input       wire                        gather_valid_i_3_22,
    output      wire                        gather_ready_o_3_22,

    output      wire        [`DW-1:0]       gather_data_o_3_22,
    output      wire                        gather_valid_o_3_22,
    input       wire                        gather_ready_i_3_22,
    input       wire        [`DW-1:0]       gather_data_i_3_23,
    input       wire                        gather_valid_i_3_23,
    output      wire                        gather_ready_o_3_23,

    output      wire        [`DW-1:0]       gather_data_o_3_23,
    output      wire                        gather_valid_o_3_23,
    input       wire                        gather_ready_i_3_23,
    input       wire        [`DW-1:0]       gather_data_i_3_24,
    input       wire                        gather_valid_i_3_24,
    output      wire                        gather_ready_o_3_24,

    output      wire        [`DW-1:0]       gather_data_o_3_24,
    output      wire                        gather_valid_o_3_24,
    input       wire                        gather_ready_i_3_24,
    input       wire        [`DW-1:0]       gather_data_i_4_0,
    input       wire                        gather_valid_i_4_0,
    output      wire                        gather_ready_o_4_0,

    output      wire        [`DW-1:0]       gather_data_o_4_0,
    output      wire                        gather_valid_o_4_0,
    input       wire                        gather_ready_i_4_0,
    input       wire        [`DW-1:0]       gather_data_i_4_1,
    input       wire                        gather_valid_i_4_1,
    output      wire                        gather_ready_o_4_1,

    output      wire        [`DW-1:0]       gather_data_o_4_1,
    output      wire                        gather_valid_o_4_1,
    input       wire                        gather_ready_i_4_1,
    input       wire        [`DW-1:0]       gather_data_i_4_2,
    input       wire                        gather_valid_i_4_2,
    output      wire                        gather_ready_o_4_2,

    output      wire        [`DW-1:0]       gather_data_o_4_2,
    output      wire                        gather_valid_o_4_2,
    input       wire                        gather_ready_i_4_2,
    input       wire        [`DW-1:0]       gather_data_i_4_3,
    input       wire                        gather_valid_i_4_3,
    output      wire                        gather_ready_o_4_3,

    output      wire        [`DW-1:0]       gather_data_o_4_3,
    output      wire                        gather_valid_o_4_3,
    input       wire                        gather_ready_i_4_3,
    input       wire        [`DW-1:0]       gather_data_i_4_4,
    input       wire                        gather_valid_i_4_4,
    output      wire                        gather_ready_o_4_4,

    output      wire        [`DW-1:0]       gather_data_o_4_4,
    output      wire                        gather_valid_o_4_4,
    input       wire                        gather_ready_i_4_4,
    input       wire        [`DW-1:0]       gather_data_i_4_5,
    input       wire                        gather_valid_i_4_5,
    output      wire                        gather_ready_o_4_5,

    output      wire        [`DW-1:0]       gather_data_o_4_5,
    output      wire                        gather_valid_o_4_5,
    input       wire                        gather_ready_i_4_5,
    input       wire        [`DW-1:0]       gather_data_i_4_6,
    input       wire                        gather_valid_i_4_6,
    output      wire                        gather_ready_o_4_6,

    output      wire        [`DW-1:0]       gather_data_o_4_6,
    output      wire                        gather_valid_o_4_6,
    input       wire                        gather_ready_i_4_6,
    input       wire        [`DW-1:0]       gather_data_i_4_7,
    input       wire                        gather_valid_i_4_7,
    output      wire                        gather_ready_o_4_7,

    output      wire        [`DW-1:0]       gather_data_o_4_7,
    output      wire                        gather_valid_o_4_7,
    input       wire                        gather_ready_i_4_7,
    input       wire        [`DW-1:0]       gather_data_i_4_8,
    input       wire                        gather_valid_i_4_8,
    output      wire                        gather_ready_o_4_8,

    output      wire        [`DW-1:0]       gather_data_o_4_8,
    output      wire                        gather_valid_o_4_8,
    input       wire                        gather_ready_i_4_8,
    input       wire        [`DW-1:0]       gather_data_i_4_9,
    input       wire                        gather_valid_i_4_9,
    output      wire                        gather_ready_o_4_9,

    output      wire        [`DW-1:0]       gather_data_o_4_9,
    output      wire                        gather_valid_o_4_9,
    input       wire                        gather_ready_i_4_9,
    input       wire        [`DW-1:0]       gather_data_i_4_10,
    input       wire                        gather_valid_i_4_10,
    output      wire                        gather_ready_o_4_10,

    output      wire        [`DW-1:0]       gather_data_o_4_10,
    output      wire                        gather_valid_o_4_10,
    input       wire                        gather_ready_i_4_10,
    input       wire        [`DW-1:0]       gather_data_i_4_11,
    input       wire                        gather_valid_i_4_11,
    output      wire                        gather_ready_o_4_11,

    output      wire        [`DW-1:0]       gather_data_o_4_11,
    output      wire                        gather_valid_o_4_11,
    input       wire                        gather_ready_i_4_11,
    input       wire        [`DW-1:0]       gather_data_i_4_12,
    input       wire                        gather_valid_i_4_12,
    output      wire                        gather_ready_o_4_12,

    output      wire        [`DW-1:0]       gather_data_o_4_12,
    output      wire                        gather_valid_o_4_12,
    input       wire                        gather_ready_i_4_12,
    input       wire        [`DW-1:0]       gather_data_i_4_13,
    input       wire                        gather_valid_i_4_13,
    output      wire                        gather_ready_o_4_13,

    output      wire        [`DW-1:0]       gather_data_o_4_13,
    output      wire                        gather_valid_o_4_13,
    input       wire                        gather_ready_i_4_13,
    input       wire        [`DW-1:0]       gather_data_i_4_14,
    input       wire                        gather_valid_i_4_14,
    output      wire                        gather_ready_o_4_14,

    output      wire        [`DW-1:0]       gather_data_o_4_14,
    output      wire                        gather_valid_o_4_14,
    input       wire                        gather_ready_i_4_14,
    input       wire        [`DW-1:0]       gather_data_i_4_15,
    input       wire                        gather_valid_i_4_15,
    output      wire                        gather_ready_o_4_15,

    output      wire        [`DW-1:0]       gather_data_o_4_15,
    output      wire                        gather_valid_o_4_15,
    input       wire                        gather_ready_i_4_15,
    input       wire        [`DW-1:0]       gather_data_i_4_16,
    input       wire                        gather_valid_i_4_16,
    output      wire                        gather_ready_o_4_16,

    output      wire        [`DW-1:0]       gather_data_o_4_16,
    output      wire                        gather_valid_o_4_16,
    input       wire                        gather_ready_i_4_16,
    input       wire        [`DW-1:0]       gather_data_i_4_17,
    input       wire                        gather_valid_i_4_17,
    output      wire                        gather_ready_o_4_17,

    output      wire        [`DW-1:0]       gather_data_o_4_17,
    output      wire                        gather_valid_o_4_17,
    input       wire                        gather_ready_i_4_17,
    input       wire        [`DW-1:0]       gather_data_i_4_18,
    input       wire                        gather_valid_i_4_18,
    output      wire                        gather_ready_o_4_18,

    output      wire        [`DW-1:0]       gather_data_o_4_18,
    output      wire                        gather_valid_o_4_18,
    input       wire                        gather_ready_i_4_18,
    input       wire        [`DW-1:0]       gather_data_i_4_19,
    input       wire                        gather_valid_i_4_19,
    output      wire                        gather_ready_o_4_19,

    output      wire        [`DW-1:0]       gather_data_o_4_19,
    output      wire                        gather_valid_o_4_19,
    input       wire                        gather_ready_i_4_19,
    input       wire        [`DW-1:0]       gather_data_i_4_20,
    input       wire                        gather_valid_i_4_20,
    output      wire                        gather_ready_o_4_20,

    output      wire        [`DW-1:0]       gather_data_o_4_20,
    output      wire                        gather_valid_o_4_20,
    input       wire                        gather_ready_i_4_20,
    input       wire        [`DW-1:0]       gather_data_i_4_21,
    input       wire                        gather_valid_i_4_21,
    output      wire                        gather_ready_o_4_21,

    output      wire        [`DW-1:0]       gather_data_o_4_21,
    output      wire                        gather_valid_o_4_21,
    input       wire                        gather_ready_i_4_21,
    input       wire        [`DW-1:0]       gather_data_i_4_22,
    input       wire                        gather_valid_i_4_22,
    output      wire                        gather_ready_o_4_22,

    output      wire        [`DW-1:0]       gather_data_o_4_22,
    output      wire                        gather_valid_o_4_22,
    input       wire                        gather_ready_i_4_22,
    input       wire        [`DW-1:0]       gather_data_i_4_23,
    input       wire                        gather_valid_i_4_23,
    output      wire                        gather_ready_o_4_23,

    output      wire        [`DW-1:0]       gather_data_o_4_23,
    output      wire                        gather_valid_o_4_23,
    input       wire                        gather_ready_i_4_23,
    input       wire        [`DW-1:0]       gather_data_i_4_24,
    input       wire                        gather_valid_i_4_24,
    output      wire                        gather_ready_o_4_24,

    output      wire        [`DW-1:0]       gather_data_o_4_24,
    output      wire                        gather_valid_o_4_24,
    input       wire                        gather_ready_i_4_24,
    input       wire        [`DW-1:0]       gather_data_i_5_0,
    input       wire                        gather_valid_i_5_0,
    output      wire                        gather_ready_o_5_0,

    output      wire        [`DW-1:0]       gather_data_o_5_0,
    output      wire                        gather_valid_o_5_0,
    input       wire                        gather_ready_i_5_0,
    input       wire        [`DW-1:0]       gather_data_i_5_1,
    input       wire                        gather_valid_i_5_1,
    output      wire                        gather_ready_o_5_1,

    output      wire        [`DW-1:0]       gather_data_o_5_1,
    output      wire                        gather_valid_o_5_1,
    input       wire                        gather_ready_i_5_1,
    input       wire        [`DW-1:0]       gather_data_i_5_2,
    input       wire                        gather_valid_i_5_2,
    output      wire                        gather_ready_o_5_2,

    output      wire        [`DW-1:0]       gather_data_o_5_2,
    output      wire                        gather_valid_o_5_2,
    input       wire                        gather_ready_i_5_2,
    input       wire        [`DW-1:0]       gather_data_i_5_3,
    input       wire                        gather_valid_i_5_3,
    output      wire                        gather_ready_o_5_3,

    output      wire        [`DW-1:0]       gather_data_o_5_3,
    output      wire                        gather_valid_o_5_3,
    input       wire                        gather_ready_i_5_3,
    input       wire        [`DW-1:0]       gather_data_i_5_4,
    input       wire                        gather_valid_i_5_4,
    output      wire                        gather_ready_o_5_4,

    output      wire        [`DW-1:0]       gather_data_o_5_4,
    output      wire                        gather_valid_o_5_4,
    input       wire                        gather_ready_i_5_4,
    input       wire        [`DW-1:0]       gather_data_i_5_5,
    input       wire                        gather_valid_i_5_5,
    output      wire                        gather_ready_o_5_5,

    output      wire        [`DW-1:0]       gather_data_o_5_5,
    output      wire                        gather_valid_o_5_5,
    input       wire                        gather_ready_i_5_5,
    input       wire        [`DW-1:0]       gather_data_i_5_6,
    input       wire                        gather_valid_i_5_6,
    output      wire                        gather_ready_o_5_6,

    output      wire        [`DW-1:0]       gather_data_o_5_6,
    output      wire                        gather_valid_o_5_6,
    input       wire                        gather_ready_i_5_6,
    input       wire        [`DW-1:0]       gather_data_i_5_7,
    input       wire                        gather_valid_i_5_7,
    output      wire                        gather_ready_o_5_7,

    output      wire        [`DW-1:0]       gather_data_o_5_7,
    output      wire                        gather_valid_o_5_7,
    input       wire                        gather_ready_i_5_7,
    input       wire        [`DW-1:0]       gather_data_i_5_8,
    input       wire                        gather_valid_i_5_8,
    output      wire                        gather_ready_o_5_8,

    output      wire        [`DW-1:0]       gather_data_o_5_8,
    output      wire                        gather_valid_o_5_8,
    input       wire                        gather_ready_i_5_8,
    input       wire        [`DW-1:0]       gather_data_i_5_9,
    input       wire                        gather_valid_i_5_9,
    output      wire                        gather_ready_o_5_9,

    output      wire        [`DW-1:0]       gather_data_o_5_9,
    output      wire                        gather_valid_o_5_9,
    input       wire                        gather_ready_i_5_9,
    input       wire        [`DW-1:0]       gather_data_i_5_10,
    input       wire                        gather_valid_i_5_10,
    output      wire                        gather_ready_o_5_10,

    output      wire        [`DW-1:0]       gather_data_o_5_10,
    output      wire                        gather_valid_o_5_10,
    input       wire                        gather_ready_i_5_10,
    input       wire        [`DW-1:0]       gather_data_i_5_11,
    input       wire                        gather_valid_i_5_11,
    output      wire                        gather_ready_o_5_11,

    output      wire        [`DW-1:0]       gather_data_o_5_11,
    output      wire                        gather_valid_o_5_11,
    input       wire                        gather_ready_i_5_11,
    input       wire        [`DW-1:0]       gather_data_i_5_12,
    input       wire                        gather_valid_i_5_12,
    output      wire                        gather_ready_o_5_12,

    output      wire        [`DW-1:0]       gather_data_o_5_12,
    output      wire                        gather_valid_o_5_12,
    input       wire                        gather_ready_i_5_12,
    input       wire        [`DW-1:0]       gather_data_i_5_13,
    input       wire                        gather_valid_i_5_13,
    output      wire                        gather_ready_o_5_13,

    output      wire        [`DW-1:0]       gather_data_o_5_13,
    output      wire                        gather_valid_o_5_13,
    input       wire                        gather_ready_i_5_13,
    input       wire        [`DW-1:0]       gather_data_i_5_14,
    input       wire                        gather_valid_i_5_14,
    output      wire                        gather_ready_o_5_14,

    output      wire        [`DW-1:0]       gather_data_o_5_14,
    output      wire                        gather_valid_o_5_14,
    input       wire                        gather_ready_i_5_14,
    input       wire        [`DW-1:0]       gather_data_i_5_15,
    input       wire                        gather_valid_i_5_15,
    output      wire                        gather_ready_o_5_15,

    output      wire        [`DW-1:0]       gather_data_o_5_15,
    output      wire                        gather_valid_o_5_15,
    input       wire                        gather_ready_i_5_15,
    input       wire        [`DW-1:0]       gather_data_i_5_16,
    input       wire                        gather_valid_i_5_16,
    output      wire                        gather_ready_o_5_16,

    output      wire        [`DW-1:0]       gather_data_o_5_16,
    output      wire                        gather_valid_o_5_16,
    input       wire                        gather_ready_i_5_16,
    input       wire        [`DW-1:0]       gather_data_i_5_17,
    input       wire                        gather_valid_i_5_17,
    output      wire                        gather_ready_o_5_17,

    output      wire        [`DW-1:0]       gather_data_o_5_17,
    output      wire                        gather_valid_o_5_17,
    input       wire                        gather_ready_i_5_17,
    input       wire        [`DW-1:0]       gather_data_i_5_18,
    input       wire                        gather_valid_i_5_18,
    output      wire                        gather_ready_o_5_18,

    output      wire        [`DW-1:0]       gather_data_o_5_18,
    output      wire                        gather_valid_o_5_18,
    input       wire                        gather_ready_i_5_18,
    input       wire        [`DW-1:0]       gather_data_i_5_19,
    input       wire                        gather_valid_i_5_19,
    output      wire                        gather_ready_o_5_19,

    output      wire        [`DW-1:0]       gather_data_o_5_19,
    output      wire                        gather_valid_o_5_19,
    input       wire                        gather_ready_i_5_19,
    input       wire        [`DW-1:0]       gather_data_i_5_20,
    input       wire                        gather_valid_i_5_20,
    output      wire                        gather_ready_o_5_20,

    output      wire        [`DW-1:0]       gather_data_o_5_20,
    output      wire                        gather_valid_o_5_20,
    input       wire                        gather_ready_i_5_20,
    input       wire        [`DW-1:0]       gather_data_i_5_21,
    input       wire                        gather_valid_i_5_21,
    output      wire                        gather_ready_o_5_21,

    output      wire        [`DW-1:0]       gather_data_o_5_21,
    output      wire                        gather_valid_o_5_21,
    input       wire                        gather_ready_i_5_21,
    input       wire        [`DW-1:0]       gather_data_i_5_22,
    input       wire                        gather_valid_i_5_22,
    output      wire                        gather_ready_o_5_22,

    output      wire        [`DW-1:0]       gather_data_o_5_22,
    output      wire                        gather_valid_o_5_22,
    input       wire                        gather_ready_i_5_22,
    input       wire        [`DW-1:0]       gather_data_i_5_23,
    input       wire                        gather_valid_i_5_23,
    output      wire                        gather_ready_o_5_23,

    output      wire        [`DW-1:0]       gather_data_o_5_23,
    output      wire                        gather_valid_o_5_23,
    input       wire                        gather_ready_i_5_23,
    input       wire        [`DW-1:0]       gather_data_i_5_24,
    input       wire                        gather_valid_i_5_24,
    output      wire                        gather_ready_o_5_24,

    output      wire        [`DW-1:0]       gather_data_o_5_24,
    output      wire                        gather_valid_o_5_24,
    input       wire                        gather_ready_i_5_24,
    input       wire        [`DW-1:0]       gather_data_i_6_0,
    input       wire                        gather_valid_i_6_0,
    output      wire                        gather_ready_o_6_0,

    output      wire        [`DW-1:0]       gather_data_o_6_0,
    output      wire                        gather_valid_o_6_0,
    input       wire                        gather_ready_i_6_0,
    input       wire        [`DW-1:0]       gather_data_i_6_1,
    input       wire                        gather_valid_i_6_1,
    output      wire                        gather_ready_o_6_1,

    output      wire        [`DW-1:0]       gather_data_o_6_1,
    output      wire                        gather_valid_o_6_1,
    input       wire                        gather_ready_i_6_1,
    input       wire        [`DW-1:0]       gather_data_i_6_2,
    input       wire                        gather_valid_i_6_2,
    output      wire                        gather_ready_o_6_2,

    output      wire        [`DW-1:0]       gather_data_o_6_2,
    output      wire                        gather_valid_o_6_2,
    input       wire                        gather_ready_i_6_2,
    input       wire        [`DW-1:0]       gather_data_i_6_3,
    input       wire                        gather_valid_i_6_3,
    output      wire                        gather_ready_o_6_3,

    output      wire        [`DW-1:0]       gather_data_o_6_3,
    output      wire                        gather_valid_o_6_3,
    input       wire                        gather_ready_i_6_3,
    input       wire        [`DW-1:0]       gather_data_i_6_4,
    input       wire                        gather_valid_i_6_4,
    output      wire                        gather_ready_o_6_4,

    output      wire        [`DW-1:0]       gather_data_o_6_4,
    output      wire                        gather_valid_o_6_4,
    input       wire                        gather_ready_i_6_4,
    input       wire        [`DW-1:0]       gather_data_i_6_5,
    input       wire                        gather_valid_i_6_5,
    output      wire                        gather_ready_o_6_5,

    output      wire        [`DW-1:0]       gather_data_o_6_5,
    output      wire                        gather_valid_o_6_5,
    input       wire                        gather_ready_i_6_5,
    input       wire        [`DW-1:0]       gather_data_i_6_6,
    input       wire                        gather_valid_i_6_6,
    output      wire                        gather_ready_o_6_6,

    output      wire        [`DW-1:0]       gather_data_o_6_6,
    output      wire                        gather_valid_o_6_6,
    input       wire                        gather_ready_i_6_6,
    input       wire        [`DW-1:0]       gather_data_i_6_7,
    input       wire                        gather_valid_i_6_7,
    output      wire                        gather_ready_o_6_7,

    output      wire        [`DW-1:0]       gather_data_o_6_7,
    output      wire                        gather_valid_o_6_7,
    input       wire                        gather_ready_i_6_7,
    input       wire        [`DW-1:0]       gather_data_i_6_8,
    input       wire                        gather_valid_i_6_8,
    output      wire                        gather_ready_o_6_8,

    output      wire        [`DW-1:0]       gather_data_o_6_8,
    output      wire                        gather_valid_o_6_8,
    input       wire                        gather_ready_i_6_8,
    input       wire        [`DW-1:0]       gather_data_i_6_9,
    input       wire                        gather_valid_i_6_9,
    output      wire                        gather_ready_o_6_9,

    output      wire        [`DW-1:0]       gather_data_o_6_9,
    output      wire                        gather_valid_o_6_9,
    input       wire                        gather_ready_i_6_9,
    input       wire        [`DW-1:0]       gather_data_i_6_10,
    input       wire                        gather_valid_i_6_10,
    output      wire                        gather_ready_o_6_10,

    output      wire        [`DW-1:0]       gather_data_o_6_10,
    output      wire                        gather_valid_o_6_10,
    input       wire                        gather_ready_i_6_10,
    input       wire        [`DW-1:0]       gather_data_i_6_11,
    input       wire                        gather_valid_i_6_11,
    output      wire                        gather_ready_o_6_11,

    output      wire        [`DW-1:0]       gather_data_o_6_11,
    output      wire                        gather_valid_o_6_11,
    input       wire                        gather_ready_i_6_11,
    input       wire        [`DW-1:0]       gather_data_i_6_12,
    input       wire                        gather_valid_i_6_12,
    output      wire                        gather_ready_o_6_12,

    output      wire        [`DW-1:0]       gather_data_o_6_12,
    output      wire                        gather_valid_o_6_12,
    input       wire                        gather_ready_i_6_12,
    input       wire        [`DW-1:0]       gather_data_i_6_13,
    input       wire                        gather_valid_i_6_13,
    output      wire                        gather_ready_o_6_13,

    output      wire        [`DW-1:0]       gather_data_o_6_13,
    output      wire                        gather_valid_o_6_13,
    input       wire                        gather_ready_i_6_13,
    input       wire        [`DW-1:0]       gather_data_i_6_14,
    input       wire                        gather_valid_i_6_14,
    output      wire                        gather_ready_o_6_14,

    output      wire        [`DW-1:0]       gather_data_o_6_14,
    output      wire                        gather_valid_o_6_14,
    input       wire                        gather_ready_i_6_14,
    input       wire        [`DW-1:0]       gather_data_i_6_15,
    input       wire                        gather_valid_i_6_15,
    output      wire                        gather_ready_o_6_15,

    output      wire        [`DW-1:0]       gather_data_o_6_15,
    output      wire                        gather_valid_o_6_15,
    input       wire                        gather_ready_i_6_15,
    input       wire        [`DW-1:0]       gather_data_i_6_16,
    input       wire                        gather_valid_i_6_16,
    output      wire                        gather_ready_o_6_16,

    output      wire        [`DW-1:0]       gather_data_o_6_16,
    output      wire                        gather_valid_o_6_16,
    input       wire                        gather_ready_i_6_16,
    input       wire        [`DW-1:0]       gather_data_i_6_17,
    input       wire                        gather_valid_i_6_17,
    output      wire                        gather_ready_o_6_17,

    output      wire        [`DW-1:0]       gather_data_o_6_17,
    output      wire                        gather_valid_o_6_17,
    input       wire                        gather_ready_i_6_17,
    input       wire        [`DW-1:0]       gather_data_i_6_18,
    input       wire                        gather_valid_i_6_18,
    output      wire                        gather_ready_o_6_18,

    output      wire        [`DW-1:0]       gather_data_o_6_18,
    output      wire                        gather_valid_o_6_18,
    input       wire                        gather_ready_i_6_18,
    input       wire        [`DW-1:0]       gather_data_i_6_19,
    input       wire                        gather_valid_i_6_19,
    output      wire                        gather_ready_o_6_19,

    output      wire        [`DW-1:0]       gather_data_o_6_19,
    output      wire                        gather_valid_o_6_19,
    input       wire                        gather_ready_i_6_19,
    input       wire        [`DW-1:0]       gather_data_i_6_20,
    input       wire                        gather_valid_i_6_20,
    output      wire                        gather_ready_o_6_20,

    output      wire        [`DW-1:0]       gather_data_o_6_20,
    output      wire                        gather_valid_o_6_20,
    input       wire                        gather_ready_i_6_20,
    input       wire        [`DW-1:0]       gather_data_i_6_21,
    input       wire                        gather_valid_i_6_21,
    output      wire                        gather_ready_o_6_21,

    output      wire        [`DW-1:0]       gather_data_o_6_21,
    output      wire                        gather_valid_o_6_21,
    input       wire                        gather_ready_i_6_21,
    input       wire        [`DW-1:0]       gather_data_i_6_22,
    input       wire                        gather_valid_i_6_22,
    output      wire                        gather_ready_o_6_22,

    output      wire        [`DW-1:0]       gather_data_o_6_22,
    output      wire                        gather_valid_o_6_22,
    input       wire                        gather_ready_i_6_22,
    input       wire        [`DW-1:0]       gather_data_i_6_23,
    input       wire                        gather_valid_i_6_23,
    output      wire                        gather_ready_o_6_23,

    output      wire        [`DW-1:0]       gather_data_o_6_23,
    output      wire                        gather_valid_o_6_23,
    input       wire                        gather_ready_i_6_23,
    input       wire        [`DW-1:0]       gather_data_i_6_24,
    input       wire                        gather_valid_i_6_24,
    output      wire                        gather_ready_o_6_24,

    output      wire        [`DW-1:0]       gather_data_o_6_24,
    output      wire                        gather_valid_o_6_24,
    input       wire                        gather_ready_i_6_24,
    input       wire        [`DW-1:0]       gather_data_i_7_0,
    input       wire                        gather_valid_i_7_0,
    output      wire                        gather_ready_o_7_0,

    output      wire        [`DW-1:0]       gather_data_o_7_0,
    output      wire                        gather_valid_o_7_0,
    input       wire                        gather_ready_i_7_0,
    input       wire        [`DW-1:0]       gather_data_i_7_1,
    input       wire                        gather_valid_i_7_1,
    output      wire                        gather_ready_o_7_1,

    output      wire        [`DW-1:0]       gather_data_o_7_1,
    output      wire                        gather_valid_o_7_1,
    input       wire                        gather_ready_i_7_1,
    input       wire        [`DW-1:0]       gather_data_i_7_2,
    input       wire                        gather_valid_i_7_2,
    output      wire                        gather_ready_o_7_2,

    output      wire        [`DW-1:0]       gather_data_o_7_2,
    output      wire                        gather_valid_o_7_2,
    input       wire                        gather_ready_i_7_2,
    input       wire        [`DW-1:0]       gather_data_i_7_3,
    input       wire                        gather_valid_i_7_3,
    output      wire                        gather_ready_o_7_3,

    output      wire        [`DW-1:0]       gather_data_o_7_3,
    output      wire                        gather_valid_o_7_3,
    input       wire                        gather_ready_i_7_3,
    input       wire        [`DW-1:0]       gather_data_i_7_4,
    input       wire                        gather_valid_i_7_4,
    output      wire                        gather_ready_o_7_4,

    output      wire        [`DW-1:0]       gather_data_o_7_4,
    output      wire                        gather_valid_o_7_4,
    input       wire                        gather_ready_i_7_4,
    input       wire        [`DW-1:0]       gather_data_i_7_5,
    input       wire                        gather_valid_i_7_5,
    output      wire                        gather_ready_o_7_5,

    output      wire        [`DW-1:0]       gather_data_o_7_5,
    output      wire                        gather_valid_o_7_5,
    input       wire                        gather_ready_i_7_5,
    input       wire        [`DW-1:0]       gather_data_i_7_6,
    input       wire                        gather_valid_i_7_6,
    output      wire                        gather_ready_o_7_6,

    output      wire        [`DW-1:0]       gather_data_o_7_6,
    output      wire                        gather_valid_o_7_6,
    input       wire                        gather_ready_i_7_6,
    input       wire        [`DW-1:0]       gather_data_i_7_7,
    input       wire                        gather_valid_i_7_7,
    output      wire                        gather_ready_o_7_7,

    output      wire        [`DW-1:0]       gather_data_o_7_7,
    output      wire                        gather_valid_o_7_7,
    input       wire                        gather_ready_i_7_7,
    input       wire        [`DW-1:0]       gather_data_i_7_8,
    input       wire                        gather_valid_i_7_8,
    output      wire                        gather_ready_o_7_8,

    output      wire        [`DW-1:0]       gather_data_o_7_8,
    output      wire                        gather_valid_o_7_8,
    input       wire                        gather_ready_i_7_8,
    input       wire        [`DW-1:0]       gather_data_i_7_9,
    input       wire                        gather_valid_i_7_9,
    output      wire                        gather_ready_o_7_9,

    output      wire        [`DW-1:0]       gather_data_o_7_9,
    output      wire                        gather_valid_o_7_9,
    input       wire                        gather_ready_i_7_9,
    input       wire        [`DW-1:0]       gather_data_i_7_10,
    input       wire                        gather_valid_i_7_10,
    output      wire                        gather_ready_o_7_10,

    output      wire        [`DW-1:0]       gather_data_o_7_10,
    output      wire                        gather_valid_o_7_10,
    input       wire                        gather_ready_i_7_10,
    input       wire        [`DW-1:0]       gather_data_i_7_11,
    input       wire                        gather_valid_i_7_11,
    output      wire                        gather_ready_o_7_11,

    output      wire        [`DW-1:0]       gather_data_o_7_11,
    output      wire                        gather_valid_o_7_11,
    input       wire                        gather_ready_i_7_11,
    input       wire        [`DW-1:0]       gather_data_i_7_12,
    input       wire                        gather_valid_i_7_12,
    output      wire                        gather_ready_o_7_12,

    output      wire        [`DW-1:0]       gather_data_o_7_12,
    output      wire                        gather_valid_o_7_12,
    input       wire                        gather_ready_i_7_12,
    input       wire        [`DW-1:0]       gather_data_i_7_13,
    input       wire                        gather_valid_i_7_13,
    output      wire                        gather_ready_o_7_13,

    output      wire        [`DW-1:0]       gather_data_o_7_13,
    output      wire                        gather_valid_o_7_13,
    input       wire                        gather_ready_i_7_13,
    input       wire        [`DW-1:0]       gather_data_i_7_14,
    input       wire                        gather_valid_i_7_14,
    output      wire                        gather_ready_o_7_14,

    output      wire        [`DW-1:0]       gather_data_o_7_14,
    output      wire                        gather_valid_o_7_14,
    input       wire                        gather_ready_i_7_14,
    input       wire        [`DW-1:0]       gather_data_i_7_15,
    input       wire                        gather_valid_i_7_15,
    output      wire                        gather_ready_o_7_15,

    output      wire        [`DW-1:0]       gather_data_o_7_15,
    output      wire                        gather_valid_o_7_15,
    input       wire                        gather_ready_i_7_15,
    input       wire        [`DW-1:0]       gather_data_i_7_16,
    input       wire                        gather_valid_i_7_16,
    output      wire                        gather_ready_o_7_16,

    output      wire        [`DW-1:0]       gather_data_o_7_16,
    output      wire                        gather_valid_o_7_16,
    input       wire                        gather_ready_i_7_16,
    input       wire        [`DW-1:0]       gather_data_i_7_17,
    input       wire                        gather_valid_i_7_17,
    output      wire                        gather_ready_o_7_17,

    output      wire        [`DW-1:0]       gather_data_o_7_17,
    output      wire                        gather_valid_o_7_17,
    input       wire                        gather_ready_i_7_17,
    input       wire        [`DW-1:0]       gather_data_i_7_18,
    input       wire                        gather_valid_i_7_18,
    output      wire                        gather_ready_o_7_18,

    output      wire        [`DW-1:0]       gather_data_o_7_18,
    output      wire                        gather_valid_o_7_18,
    input       wire                        gather_ready_i_7_18,
    input       wire        [`DW-1:0]       gather_data_i_7_19,
    input       wire                        gather_valid_i_7_19,
    output      wire                        gather_ready_o_7_19,

    output      wire        [`DW-1:0]       gather_data_o_7_19,
    output      wire                        gather_valid_o_7_19,
    input       wire                        gather_ready_i_7_19,
    input       wire        [`DW-1:0]       gather_data_i_7_20,
    input       wire                        gather_valid_i_7_20,
    output      wire                        gather_ready_o_7_20,

    output      wire        [`DW-1:0]       gather_data_o_7_20,
    output      wire                        gather_valid_o_7_20,
    input       wire                        gather_ready_i_7_20,
    input       wire        [`DW-1:0]       gather_data_i_7_21,
    input       wire                        gather_valid_i_7_21,
    output      wire                        gather_ready_o_7_21,

    output      wire        [`DW-1:0]       gather_data_o_7_21,
    output      wire                        gather_valid_o_7_21,
    input       wire                        gather_ready_i_7_21,
    input       wire        [`DW-1:0]       gather_data_i_7_22,
    input       wire                        gather_valid_i_7_22,
    output      wire                        gather_ready_o_7_22,

    output      wire        [`DW-1:0]       gather_data_o_7_22,
    output      wire                        gather_valid_o_7_22,
    input       wire                        gather_ready_i_7_22,
    input       wire        [`DW-1:0]       gather_data_i_7_23,
    input       wire                        gather_valid_i_7_23,
    output      wire                        gather_ready_o_7_23,

    output      wire        [`DW-1:0]       gather_data_o_7_23,
    output      wire                        gather_valid_o_7_23,
    input       wire                        gather_ready_i_7_23,
    input       wire        [`DW-1:0]       gather_data_i_7_24,
    input       wire                        gather_valid_i_7_24,
    output      wire                        gather_ready_o_7_24,

    output      wire        [`DW-1:0]       gather_data_o_7_24,
    output      wire                        gather_valid_o_7_24,
    input       wire                        gather_ready_i_7_24,
    input       wire        [`DW-1:0]       gather_data_i_8_0,
    input       wire                        gather_valid_i_8_0,
    output      wire                        gather_ready_o_8_0,

    output      wire        [`DW-1:0]       gather_data_o_8_0,
    output      wire                        gather_valid_o_8_0,
    input       wire                        gather_ready_i_8_0,
    input       wire        [`DW-1:0]       gather_data_i_8_1,
    input       wire                        gather_valid_i_8_1,
    output      wire                        gather_ready_o_8_1,

    output      wire        [`DW-1:0]       gather_data_o_8_1,
    output      wire                        gather_valid_o_8_1,
    input       wire                        gather_ready_i_8_1,
    input       wire        [`DW-1:0]       gather_data_i_8_2,
    input       wire                        gather_valid_i_8_2,
    output      wire                        gather_ready_o_8_2,

    output      wire        [`DW-1:0]       gather_data_o_8_2,
    output      wire                        gather_valid_o_8_2,
    input       wire                        gather_ready_i_8_2,
    input       wire        [`DW-1:0]       gather_data_i_8_3,
    input       wire                        gather_valid_i_8_3,
    output      wire                        gather_ready_o_8_3,

    output      wire        [`DW-1:0]       gather_data_o_8_3,
    output      wire                        gather_valid_o_8_3,
    input       wire                        gather_ready_i_8_3,
    input       wire        [`DW-1:0]       gather_data_i_8_4,
    input       wire                        gather_valid_i_8_4,
    output      wire                        gather_ready_o_8_4,

    output      wire        [`DW-1:0]       gather_data_o_8_4,
    output      wire                        gather_valid_o_8_4,
    input       wire                        gather_ready_i_8_4,
    input       wire        [`DW-1:0]       gather_data_i_8_5,
    input       wire                        gather_valid_i_8_5,
    output      wire                        gather_ready_o_8_5,

    output      wire        [`DW-1:0]       gather_data_o_8_5,
    output      wire                        gather_valid_o_8_5,
    input       wire                        gather_ready_i_8_5,
    input       wire        [`DW-1:0]       gather_data_i_8_6,
    input       wire                        gather_valid_i_8_6,
    output      wire                        gather_ready_o_8_6,

    output      wire        [`DW-1:0]       gather_data_o_8_6,
    output      wire                        gather_valid_o_8_6,
    input       wire                        gather_ready_i_8_6,
    input       wire        [`DW-1:0]       gather_data_i_8_7,
    input       wire                        gather_valid_i_8_7,
    output      wire                        gather_ready_o_8_7,

    output      wire        [`DW-1:0]       gather_data_o_8_7,
    output      wire                        gather_valid_o_8_7,
    input       wire                        gather_ready_i_8_7,
    input       wire        [`DW-1:0]       gather_data_i_8_8,
    input       wire                        gather_valid_i_8_8,
    output      wire                        gather_ready_o_8_8,

    output      wire        [`DW-1:0]       gather_data_o_8_8,
    output      wire                        gather_valid_o_8_8,
    input       wire                        gather_ready_i_8_8,
    input       wire        [`DW-1:0]       gather_data_i_8_9,
    input       wire                        gather_valid_i_8_9,
    output      wire                        gather_ready_o_8_9,

    output      wire        [`DW-1:0]       gather_data_o_8_9,
    output      wire                        gather_valid_o_8_9,
    input       wire                        gather_ready_i_8_9,
    input       wire        [`DW-1:0]       gather_data_i_8_10,
    input       wire                        gather_valid_i_8_10,
    output      wire                        gather_ready_o_8_10,

    output      wire        [`DW-1:0]       gather_data_o_8_10,
    output      wire                        gather_valid_o_8_10,
    input       wire                        gather_ready_i_8_10,
    input       wire        [`DW-1:0]       gather_data_i_8_11,
    input       wire                        gather_valid_i_8_11,
    output      wire                        gather_ready_o_8_11,

    output      wire        [`DW-1:0]       gather_data_o_8_11,
    output      wire                        gather_valid_o_8_11,
    input       wire                        gather_ready_i_8_11,
    input       wire        [`DW-1:0]       gather_data_i_8_12,
    input       wire                        gather_valid_i_8_12,
    output      wire                        gather_ready_o_8_12,

    output      wire        [`DW-1:0]       gather_data_o_8_12,
    output      wire                        gather_valid_o_8_12,
    input       wire                        gather_ready_i_8_12,
    input       wire        [`DW-1:0]       gather_data_i_8_13,
    input       wire                        gather_valid_i_8_13,
    output      wire                        gather_ready_o_8_13,

    output      wire        [`DW-1:0]       gather_data_o_8_13,
    output      wire                        gather_valid_o_8_13,
    input       wire                        gather_ready_i_8_13,
    input       wire        [`DW-1:0]       gather_data_i_8_14,
    input       wire                        gather_valid_i_8_14,
    output      wire                        gather_ready_o_8_14,

    output      wire        [`DW-1:0]       gather_data_o_8_14,
    output      wire                        gather_valid_o_8_14,
    input       wire                        gather_ready_i_8_14,
    input       wire        [`DW-1:0]       gather_data_i_8_15,
    input       wire                        gather_valid_i_8_15,
    output      wire                        gather_ready_o_8_15,

    output      wire        [`DW-1:0]       gather_data_o_8_15,
    output      wire                        gather_valid_o_8_15,
    input       wire                        gather_ready_i_8_15,
    input       wire        [`DW-1:0]       gather_data_i_8_16,
    input       wire                        gather_valid_i_8_16,
    output      wire                        gather_ready_o_8_16,

    output      wire        [`DW-1:0]       gather_data_o_8_16,
    output      wire                        gather_valid_o_8_16,
    input       wire                        gather_ready_i_8_16,
    input       wire        [`DW-1:0]       gather_data_i_8_17,
    input       wire                        gather_valid_i_8_17,
    output      wire                        gather_ready_o_8_17,

    output      wire        [`DW-1:0]       gather_data_o_8_17,
    output      wire                        gather_valid_o_8_17,
    input       wire                        gather_ready_i_8_17,
    input       wire        [`DW-1:0]       gather_data_i_8_18,
    input       wire                        gather_valid_i_8_18,
    output      wire                        gather_ready_o_8_18,

    output      wire        [`DW-1:0]       gather_data_o_8_18,
    output      wire                        gather_valid_o_8_18,
    input       wire                        gather_ready_i_8_18,
    input       wire        [`DW-1:0]       gather_data_i_8_19,
    input       wire                        gather_valid_i_8_19,
    output      wire                        gather_ready_o_8_19,

    output      wire        [`DW-1:0]       gather_data_o_8_19,
    output      wire                        gather_valid_o_8_19,
    input       wire                        gather_ready_i_8_19,
    input       wire        [`DW-1:0]       gather_data_i_8_20,
    input       wire                        gather_valid_i_8_20,
    output      wire                        gather_ready_o_8_20,

    output      wire        [`DW-1:0]       gather_data_o_8_20,
    output      wire                        gather_valid_o_8_20,
    input       wire                        gather_ready_i_8_20,
    input       wire        [`DW-1:0]       gather_data_i_8_21,
    input       wire                        gather_valid_i_8_21,
    output      wire                        gather_ready_o_8_21,

    output      wire        [`DW-1:0]       gather_data_o_8_21,
    output      wire                        gather_valid_o_8_21,
    input       wire                        gather_ready_i_8_21,
    input       wire        [`DW-1:0]       gather_data_i_8_22,
    input       wire                        gather_valid_i_8_22,
    output      wire                        gather_ready_o_8_22,

    output      wire        [`DW-1:0]       gather_data_o_8_22,
    output      wire                        gather_valid_o_8_22,
    input       wire                        gather_ready_i_8_22,
    input       wire        [`DW-1:0]       gather_data_i_8_23,
    input       wire                        gather_valid_i_8_23,
    output      wire                        gather_ready_o_8_23,

    output      wire        [`DW-1:0]       gather_data_o_8_23,
    output      wire                        gather_valid_o_8_23,
    input       wire                        gather_ready_i_8_23,
    input       wire        [`DW-1:0]       gather_data_i_8_24,
    input       wire                        gather_valid_i_8_24,
    output      wire                        gather_ready_o_8_24,

    output      wire        [`DW-1:0]       gather_data_o_8_24,
    output      wire                        gather_valid_o_8_24,
    input       wire                        gather_ready_i_8_24,
    input       wire        [`DW-1:0]       gather_data_i_9_0,
    input       wire                        gather_valid_i_9_0,
    output      wire                        gather_ready_o_9_0,

    output      wire        [`DW-1:0]       gather_data_o_9_0,
    output      wire                        gather_valid_o_9_0,
    input       wire                        gather_ready_i_9_0,
    input       wire        [`DW-1:0]       gather_data_i_9_1,
    input       wire                        gather_valid_i_9_1,
    output      wire                        gather_ready_o_9_1,

    output      wire        [`DW-1:0]       gather_data_o_9_1,
    output      wire                        gather_valid_o_9_1,
    input       wire                        gather_ready_i_9_1,
    input       wire        [`DW-1:0]       gather_data_i_9_2,
    input       wire                        gather_valid_i_9_2,
    output      wire                        gather_ready_o_9_2,

    output      wire        [`DW-1:0]       gather_data_o_9_2,
    output      wire                        gather_valid_o_9_2,
    input       wire                        gather_ready_i_9_2,
    input       wire        [`DW-1:0]       gather_data_i_9_3,
    input       wire                        gather_valid_i_9_3,
    output      wire                        gather_ready_o_9_3,

    output      wire        [`DW-1:0]       gather_data_o_9_3,
    output      wire                        gather_valid_o_9_3,
    input       wire                        gather_ready_i_9_3,
    input       wire        [`DW-1:0]       gather_data_i_9_4,
    input       wire                        gather_valid_i_9_4,
    output      wire                        gather_ready_o_9_4,

    output      wire        [`DW-1:0]       gather_data_o_9_4,
    output      wire                        gather_valid_o_9_4,
    input       wire                        gather_ready_i_9_4,
    input       wire        [`DW-1:0]       gather_data_i_9_5,
    input       wire                        gather_valid_i_9_5,
    output      wire                        gather_ready_o_9_5,

    output      wire        [`DW-1:0]       gather_data_o_9_5,
    output      wire                        gather_valid_o_9_5,
    input       wire                        gather_ready_i_9_5,
    input       wire        [`DW-1:0]       gather_data_i_9_6,
    input       wire                        gather_valid_i_9_6,
    output      wire                        gather_ready_o_9_6,

    output      wire        [`DW-1:0]       gather_data_o_9_6,
    output      wire                        gather_valid_o_9_6,
    input       wire                        gather_ready_i_9_6,
    input       wire        [`DW-1:0]       gather_data_i_9_7,
    input       wire                        gather_valid_i_9_7,
    output      wire                        gather_ready_o_9_7,

    output      wire        [`DW-1:0]       gather_data_o_9_7,
    output      wire                        gather_valid_o_9_7,
    input       wire                        gather_ready_i_9_7,
    input       wire        [`DW-1:0]       gather_data_i_9_8,
    input       wire                        gather_valid_i_9_8,
    output      wire                        gather_ready_o_9_8,

    output      wire        [`DW-1:0]       gather_data_o_9_8,
    output      wire                        gather_valid_o_9_8,
    input       wire                        gather_ready_i_9_8,
    input       wire        [`DW-1:0]       gather_data_i_9_9,
    input       wire                        gather_valid_i_9_9,
    output      wire                        gather_ready_o_9_9,

    output      wire        [`DW-1:0]       gather_data_o_9_9,
    output      wire                        gather_valid_o_9_9,
    input       wire                        gather_ready_i_9_9,
    input       wire        [`DW-1:0]       gather_data_i_9_10,
    input       wire                        gather_valid_i_9_10,
    output      wire                        gather_ready_o_9_10,

    output      wire        [`DW-1:0]       gather_data_o_9_10,
    output      wire                        gather_valid_o_9_10,
    input       wire                        gather_ready_i_9_10,
    input       wire        [`DW-1:0]       gather_data_i_9_11,
    input       wire                        gather_valid_i_9_11,
    output      wire                        gather_ready_o_9_11,

    output      wire        [`DW-1:0]       gather_data_o_9_11,
    output      wire                        gather_valid_o_9_11,
    input       wire                        gather_ready_i_9_11,
    input       wire        [`DW-1:0]       gather_data_i_9_12,
    input       wire                        gather_valid_i_9_12,
    output      wire                        gather_ready_o_9_12,

    output      wire        [`DW-1:0]       gather_data_o_9_12,
    output      wire                        gather_valid_o_9_12,
    input       wire                        gather_ready_i_9_12,
    input       wire        [`DW-1:0]       gather_data_i_9_13,
    input       wire                        gather_valid_i_9_13,
    output      wire                        gather_ready_o_9_13,

    output      wire        [`DW-1:0]       gather_data_o_9_13,
    output      wire                        gather_valid_o_9_13,
    input       wire                        gather_ready_i_9_13,
    input       wire        [`DW-1:0]       gather_data_i_9_14,
    input       wire                        gather_valid_i_9_14,
    output      wire                        gather_ready_o_9_14,

    output      wire        [`DW-1:0]       gather_data_o_9_14,
    output      wire                        gather_valid_o_9_14,
    input       wire                        gather_ready_i_9_14,
    input       wire        [`DW-1:0]       gather_data_i_9_15,
    input       wire                        gather_valid_i_9_15,
    output      wire                        gather_ready_o_9_15,

    output      wire        [`DW-1:0]       gather_data_o_9_15,
    output      wire                        gather_valid_o_9_15,
    input       wire                        gather_ready_i_9_15,
    input       wire        [`DW-1:0]       gather_data_i_9_16,
    input       wire                        gather_valid_i_9_16,
    output      wire                        gather_ready_o_9_16,

    output      wire        [`DW-1:0]       gather_data_o_9_16,
    output      wire                        gather_valid_o_9_16,
    input       wire                        gather_ready_i_9_16,
    input       wire        [`DW-1:0]       gather_data_i_9_17,
    input       wire                        gather_valid_i_9_17,
    output      wire                        gather_ready_o_9_17,

    output      wire        [`DW-1:0]       gather_data_o_9_17,
    output      wire                        gather_valid_o_9_17,
    input       wire                        gather_ready_i_9_17,
    input       wire        [`DW-1:0]       gather_data_i_9_18,
    input       wire                        gather_valid_i_9_18,
    output      wire                        gather_ready_o_9_18,

    output      wire        [`DW-1:0]       gather_data_o_9_18,
    output      wire                        gather_valid_o_9_18,
    input       wire                        gather_ready_i_9_18,
    input       wire        [`DW-1:0]       gather_data_i_9_19,
    input       wire                        gather_valid_i_9_19,
    output      wire                        gather_ready_o_9_19,

    output      wire        [`DW-1:0]       gather_data_o_9_19,
    output      wire                        gather_valid_o_9_19,
    input       wire                        gather_ready_i_9_19,
    input       wire        [`DW-1:0]       gather_data_i_9_20,
    input       wire                        gather_valid_i_9_20,
    output      wire                        gather_ready_o_9_20,

    output      wire        [`DW-1:0]       gather_data_o_9_20,
    output      wire                        gather_valid_o_9_20,
    input       wire                        gather_ready_i_9_20,
    input       wire        [`DW-1:0]       gather_data_i_9_21,
    input       wire                        gather_valid_i_9_21,
    output      wire                        gather_ready_o_9_21,

    output      wire        [`DW-1:0]       gather_data_o_9_21,
    output      wire                        gather_valid_o_9_21,
    input       wire                        gather_ready_i_9_21,
    input       wire        [`DW-1:0]       gather_data_i_9_22,
    input       wire                        gather_valid_i_9_22,
    output      wire                        gather_ready_o_9_22,

    output      wire        [`DW-1:0]       gather_data_o_9_22,
    output      wire                        gather_valid_o_9_22,
    input       wire                        gather_ready_i_9_22,
    input       wire        [`DW-1:0]       gather_data_i_9_23,
    input       wire                        gather_valid_i_9_23,
    output      wire                        gather_ready_o_9_23,

    output      wire        [`DW-1:0]       gather_data_o_9_23,
    output      wire                        gather_valid_o_9_23,
    input       wire                        gather_ready_i_9_23,
    input       wire        [`DW-1:0]       gather_data_i_9_24,
    input       wire                        gather_valid_i_9_24,
    output      wire                        gather_ready_o_9_24,

    output      wire        [`DW-1:0]       gather_data_o_9_24,
    output      wire                        gather_valid_o_9_24,
    input       wire                        gather_ready_i_9_24
);
wire [`DW-1:0] data_stab;
wire valid_stab, ready_stab;

wire [`DW-1:0] data_flee0;
wire valid_flee0, ready_flee0;

wire [`DW-1:0] data_flee1;
wire valid_flee1, ready_flee1;

wire [`DW-1:0] data_flee2;
wire valid_flee2, ready_flee2;

wire [`DW-1:0] data_flee3;
wire valid_flee3, ready_flee3;

wire [`DW-1:0] data_flee4;
wire valid_flee4, ready_flee4;

wire [`DW-1:0] data_flee5;
wire valid_flee5, ready_flee5;

wire [`DW-1:0] data_flee6;
wire valid_flee6, ready_flee6;

wire [`DW-1:0] data_flee7;
wire valid_flee7, ready_flee7;

wire [`DW-1:0] data_i_cast_nw[`NOC_WIDTH][`NOC_HEIGHT], data_o_cast_nw[`NOC_WIDTH][`NOC_HEIGHT], data_i_merge_nw[`NOC_WIDTH][`NOC_HEIGHT], data_o_merge_nw[`NOC_WIDTH][`NOC_HEIGHT], data_i_gather_nw[`NOC_WIDTH][`NOC_HEIGHT], data_o_gather_nw[`NOC_WIDTH][`NOC_HEIGHT];
wire valid_i_cast_nw[`NOC_WIDTH][`NOC_HEIGHT], valid_o_cast_nw[`NOC_WIDTH][`NOC_HEIGHT], valid_i_merge_nw[`NOC_WIDTH][`NOC_HEIGHT], valid_o_merge_nw[`NOC_WIDTH][`NOC_HEIGHT], valid_i_gather_nw[`NOC_WIDTH][`NOC_HEIGHT], valid_o_gather_nw[`NOC_WIDTH][`NOC_HEIGHT];
wire ready_i_cast_nw[`NOC_WIDTH][`NOC_HEIGHT], ready_o_cast_nw[`NOC_WIDTH][`NOC_HEIGHT], ready_i_merge_nw[`NOC_WIDTH][`NOC_HEIGHT], ready_o_merge_nw[`NOC_WIDTH][`NOC_HEIGHT], ready_i_gather_nw[`NOC_WIDTH][`NOC_HEIGHT], ready_o_gather_nw[`NOC_WIDTH][`NOC_HEIGHT];

wire credit_upd[`NOC_WIDTH][`NOC_HEIGHT];

// from stab port to network
converter #(
    .out                            (1),
    .sid                            (1023)
)converter_stab(
    .clk                            (clk),
    .rstn                           (rstn),
    .valid_i_pe                     (valid_i_stab),
    .data_i_pe                      (data_i_stab),
    .ready_o_pe                     (ready_o_stab),
    .valid_o_pe                     (),
    .data_o_pe                      (),
    .ready_i_pe                     (1'b0),
    .valid_i_nw                     (1'b0),
    .data_i_nw                      ({(`DW){1'b0}}),
    .ready_o_nw                     (),
    .valid_o_nw                     (valid_stab),
    .data_o_nw                      (data_stab),
    .ready_i_nw                     (ready_stab)
);

// from flee0 port to outside
converter #(
    .out                            (0),
    .sid                            (1022)
)converter_flee0(
    .clk                            (clk),
    .rstn                           (rstn),
    .valid_i_pe                     (1'b0),
    .data_i_pe                      ({(`DW){1'b0}}),
    .ready_o_pe                     (),
    .valid_o_pe                     (valid_o_flee0),
    .data_o_pe                      (data_o_flee0),
    .ready_i_pe                     (ready_i_flee0),
    .valid_i_nw                     (valid_flee0),
    .data_i_nw                      (data_flee0),
    .ready_o_nw                     (ready_flee0),
    .valid_o_nw                     (),
    .data_o_nw                      (),
    .ready_i_nw                     (1'b0)
);

// from flee1 port to outside
converter #(
    .out                            (0),
    .sid                            (1022)
)converter_flee1(
    .clk                            (clk),
    .rstn                           (rstn),
    .valid_i_pe                     (1'b0),
    .data_i_pe                      ({(`DW){1'b0}}),
    .ready_o_pe                     (),
    .valid_o_pe                     (valid_o_flee1),
    .data_o_pe                      (data_o_flee1),
    .ready_i_pe                     (ready_i_flee1),
    .valid_i_nw                     (valid_flee1),
    .data_i_nw                      (data_flee1),
    .ready_o_nw                     (ready_flee1),
    .valid_o_nw                     (),
    .data_o_nw                      (),
    .ready_i_nw                     (1'b0)
);

// from flee2 port to outside
converter #(
    .out                            (0),
    .sid                            (1022)
)converter_flee2(
    .clk                            (clk),
    .rstn                           (rstn),
    .valid_i_pe                     (1'b0),
    .data_i_pe                      ({(`DW){1'b0}}),
    .ready_o_pe                     (),
    .valid_o_pe                     (valid_o_flee2),
    .data_o_pe                      (data_o_flee2),
    .ready_i_pe                     (ready_i_flee2),
    .valid_i_nw                     (valid_flee2),
    .data_i_nw                      (data_flee2),
    .ready_o_nw                     (ready_flee2),
    .valid_o_nw                     (),
    .data_o_nw                      (),
    .ready_i_nw                     (1'b0)
);

// from flee3 port to outside
converter #(
    .out                            (0),
    .sid                            (1022)
)converter_flee3(
    .clk                            (clk),
    .rstn                           (rstn),
    .valid_i_pe                     (1'b0),
    .data_i_pe                      ({(`DW){1'b0}}),
    .ready_o_pe                     (),
    .valid_o_pe                     (valid_o_flee3),
    .data_o_pe                      (data_o_flee3),
    .ready_i_pe                     (ready_i_flee3),
    .valid_i_nw                     (valid_flee3),
    .data_i_nw                      (data_flee3),
    .ready_o_nw                     (ready_flee3),
    .valid_o_nw                     (),
    .data_o_nw                      (),
    .ready_i_nw                     (1'b0)
);

// from flee4 port to outside
converter #(
    .out                            (0),
    .sid                            (1022)
)converter_flee4(
    .clk                            (clk),
    .rstn                           (rstn),
    .valid_i_pe                     (1'b0),
    .data_i_pe                      ({(`DW){1'b0}}),
    .ready_o_pe                     (),
    .valid_o_pe                     (valid_o_flee4),
    .data_o_pe                      (data_o_flee4),
    .ready_i_pe                     (ready_i_flee4),
    .valid_i_nw                     (valid_flee4),
    .data_i_nw                      (data_flee4),
    .ready_o_nw                     (ready_flee4),
    .valid_o_nw                     (),
    .data_o_nw                      (),
    .ready_i_nw                     (1'b0)
);

// from flee5 port to outside
converter #(
    .out                            (0),
    .sid                            (1022)
)converter_flee5(
    .clk                            (clk),
    .rstn                           (rstn),
    .valid_i_pe                     (1'b0),
    .data_i_pe                      ({(`DW){1'b0}}),
    .ready_o_pe                     (),
    .valid_o_pe                     (valid_o_flee5),
    .data_o_pe                      (data_o_flee5),
    .ready_i_pe                     (ready_i_flee5),
    .valid_i_nw                     (valid_flee5),
    .data_i_nw                      (data_flee5),
    .ready_o_nw                     (ready_flee5),
    .valid_o_nw                     (),
    .data_o_nw                      (),
    .ready_i_nw                     (1'b0)
);

// from flee6 port to outside
converter #(
    .out                            (0),
    .sid                            (1022)
)converter_flee6(
    .clk                            (clk),
    .rstn                           (rstn),
    .valid_i_pe                     (1'b0),
    .data_i_pe                      ({(`DW){1'b0}}),
    .ready_o_pe                     (),
    .valid_o_pe                     (valid_o_flee6),
    .data_o_pe                      (data_o_flee6),
    .ready_i_pe                     (ready_i_flee6),
    .valid_i_nw                     (valid_flee6),
    .data_i_nw                      (data_flee6),
    .ready_o_nw                     (ready_flee6),
    .valid_o_nw                     (),
    .data_o_nw                      (),
    .ready_i_nw                     (1'b0)
);

// from flee7 port to outside
converter #(
    .out                            (0),
    .sid                            (1022)
)converter_flee7(
    .clk                            (clk),
    .rstn                           (rstn),
    .valid_i_pe                     (1'b0),
    .data_i_pe                      ({(`DW){1'b0}}),
    .ready_o_pe                     (),
    .valid_o_pe                     (valid_o_flee7),
    .data_o_pe                      (data_o_flee7),
    .ready_i_pe                     (ready_i_flee7),
    .valid_i_nw                     (valid_flee7),
    .data_i_nw                      (data_flee7),
    .ready_o_nw                     (ready_flee7),
    .valid_o_nw                     (),
    .data_o_nw                      (),
    .ready_i_nw                     (1'b0)
);

cast_network cast_nw(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_cast_nw),
    .valid_i                        (valid_i_cast_nw),
    .ready_o                        (ready_o_cast_nw),
    .data_o                         (data_o_cast_nw),
    .valid_o                        (valid_o_cast_nw),
    .ready_i                        (ready_i_cast_nw),
    .data_i_stab                    (data_stab),
    .valid_i_stab                   (valid_stab),
    .ready_o_stab                   (ready_stab),
    .data_o_flee0                   (data_flee0),
    .valid_o_flee0                  (valid_flee0),
    .ready_i_flee0                  (ready_flee0),
    .data_o_flee1                   (data_flee1),
    .valid_o_flee1                  (valid_flee1),
    .ready_i_flee1                  (ready_flee1),
    .data_o_flee2                   (data_flee2),
    .valid_o_flee2                  (valid_flee2),
    .ready_i_flee2                  (ready_flee2),
    .data_o_flee3                   (data_flee3),
    .valid_o_flee3                  (valid_flee3),
    .ready_i_flee3                  (ready_flee3),
    .data_o_flee4                   (data_flee4),
    .valid_o_flee4                  (valid_flee4),
    .ready_i_flee4                  (ready_flee4),
    .data_o_flee5                   (data_flee5),
    .valid_o_flee5                  (valid_flee5),
    .ready_i_flee5                  (ready_flee5),
    .data_o_flee6                   (data_flee6),
    .valid_o_flee6                  (valid_flee6),
    .ready_i_flee6                  (ready_flee6),
    .data_o_flee7                   (data_flee7),
    .valid_o_flee7                  (valid_flee7),
    .ready_i_flee7                  (ready_flee7),
    .credit_upd                     (credit_upd)
);                 

merge_network merge_nw(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_merge_nw),
    .valid_i                        (valid_i_merge_nw),
    .ready_o                        (ready_o_merge_nw),
    .data_o                         (data_o_merge_nw),
    .valid_o                        (valid_o_merge_nw),
    .ready_i                        (ready_i_merge_nw)
);

gather_network gather_nw(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_gather_nw),
    .valid_i                        (valid_i_gather_nw),
    .ready_o                        (ready_o_gather_nw),
    .data_o                         (data_o_gather_nw),
    .valid_o                        (valid_o_gather_nw),
    .ready_i                        (ready_i_gather_nw)
);


network_interface #(
    .cast_out                       (cast_out_0_0),
    .gather_out                     (gather_out_0_0),
    .cast_sid                       (cast_sid_0_0),
    .gather_sid                     (gather_sid_0_0)
)ni_0_0(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[0][0]),
    .data_i_cast_nw                 (data_o_cast_nw[0][0]),
    .ready_o_cast_nw                (ready_i_cast_nw[0][0]),
    .valid_o_cast_nw                (valid_i_cast_nw[0][0]),
    .data_o_cast_nw                 (data_i_cast_nw[0][0]),
    .ready_i_cast_nw                (ready_o_cast_nw[0][0]),

    .valid_i_gather_nw              (valid_o_gather_nw[0][0]),
    .data_i_gather_nw               (data_o_gather_nw[0][0]),
    .ready_o_gather_nw              (ready_i_gather_nw[0][0]),
    .valid_o_gather_nw              (valid_i_gather_nw[0][0]),
    .data_o_gather_nw               (data_i_gather_nw[0][0]),
    .ready_i_gather_nw              (ready_o_gather_nw[0][0]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[0][0]),
    .data_i_merge_nw                (data_o_merge_nw[0][0]),
    .ready_o_merge_nw               (ready_i_merge_nw[0][0]),
    .valid_o_merge_nw               (valid_i_merge_nw[0][0]),
    .data_o_merge_nw                (data_i_merge_nw[0][0]),
    .ready_i_merge_nw               (ready_o_merge_nw[0][0]),

    .valid_i_cast_pe                (cast_valid_i_0_0),
    .data_i_cast_pe                 (cast_data_i_0_0),
    .ready_o_cast_pe                (cast_ready_o_0_0),
    .valid_o_cast_pe                (cast_valid_o_0_0),
    .data_o_cast_pe                 (cast_data_o_0_0),
    .ready_i_cast_pe                (cast_ready_i_0_0),

    .valid_i_merge_pe               (merge_valid_i_0_0),
    .data_i_merge_pe                (merge_data_i_0_0),
    .ready_o_merge_pe               (merge_ready_o_0_0),
    .valid_o_merge_pe               (merge_valid_o_0_0),
    .data_o_merge_pe                (merge_data_o_0_0),
    .ready_i_merge_pe               (merge_ready_i_0_0),

    .valid_i_gather_pe              (gather_valid_i_0_0),
    .data_i_gather_pe               (gather_data_i_0_0),
    .ready_o_gather_pe              (gather_ready_o_0_0),
    .valid_o_gather_pe              (gather_valid_o_0_0),
    .data_o_gather_pe               (gather_data_o_0_0),
    .ready_i_gather_pe              (gather_ready_i_0_0),

    .credit_upd                     (credit_upd[0][0])
);


network_interface #(
    .cast_out                       (cast_out_0_1),
    .gather_out                     (gather_out_0_1),
    .cast_sid                       (cast_sid_0_1),
    .gather_sid                     (gather_sid_0_1)
)ni_0_1(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[0][1]),
    .data_i_cast_nw                 (data_o_cast_nw[0][1]),
    .ready_o_cast_nw                (ready_i_cast_nw[0][1]),
    .valid_o_cast_nw                (valid_i_cast_nw[0][1]),
    .data_o_cast_nw                 (data_i_cast_nw[0][1]),
    .ready_i_cast_nw                (ready_o_cast_nw[0][1]),

    .valid_i_gather_nw              (valid_o_gather_nw[0][1]),
    .data_i_gather_nw               (data_o_gather_nw[0][1]),
    .ready_o_gather_nw              (ready_i_gather_nw[0][1]),
    .valid_o_gather_nw              (valid_i_gather_nw[0][1]),
    .data_o_gather_nw               (data_i_gather_nw[0][1]),
    .ready_i_gather_nw              (ready_o_gather_nw[0][1]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[0][1]),
    .data_i_merge_nw                (data_o_merge_nw[0][1]),
    .ready_o_merge_nw               (ready_i_merge_nw[0][1]),
    .valid_o_merge_nw               (valid_i_merge_nw[0][1]),
    .data_o_merge_nw                (data_i_merge_nw[0][1]),
    .ready_i_merge_nw               (ready_o_merge_nw[0][1]),

    .valid_i_cast_pe                (cast_valid_i_0_1),
    .data_i_cast_pe                 (cast_data_i_0_1),
    .ready_o_cast_pe                (cast_ready_o_0_1),
    .valid_o_cast_pe                (cast_valid_o_0_1),
    .data_o_cast_pe                 (cast_data_o_0_1),
    .ready_i_cast_pe                (cast_ready_i_0_1),

    .valid_i_merge_pe               (merge_valid_i_0_1),
    .data_i_merge_pe                (merge_data_i_0_1),
    .ready_o_merge_pe               (merge_ready_o_0_1),
    .valid_o_merge_pe               (merge_valid_o_0_1),
    .data_o_merge_pe                (merge_data_o_0_1),
    .ready_i_merge_pe               (merge_ready_i_0_1),

    .valid_i_gather_pe              (gather_valid_i_0_1),
    .data_i_gather_pe               (gather_data_i_0_1),
    .ready_o_gather_pe              (gather_ready_o_0_1),
    .valid_o_gather_pe              (gather_valid_o_0_1),
    .data_o_gather_pe               (gather_data_o_0_1),
    .ready_i_gather_pe              (gather_ready_i_0_1),

    .credit_upd                     (credit_upd[0][1])
);


network_interface #(
    .cast_out                       (cast_out_0_2),
    .gather_out                     (gather_out_0_2),
    .cast_sid                       (cast_sid_0_2),
    .gather_sid                     (gather_sid_0_2)
)ni_0_2(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[0][2]),
    .data_i_cast_nw                 (data_o_cast_nw[0][2]),
    .ready_o_cast_nw                (ready_i_cast_nw[0][2]),
    .valid_o_cast_nw                (valid_i_cast_nw[0][2]),
    .data_o_cast_nw                 (data_i_cast_nw[0][2]),
    .ready_i_cast_nw                (ready_o_cast_nw[0][2]),

    .valid_i_gather_nw              (valid_o_gather_nw[0][2]),
    .data_i_gather_nw               (data_o_gather_nw[0][2]),
    .ready_o_gather_nw              (ready_i_gather_nw[0][2]),
    .valid_o_gather_nw              (valid_i_gather_nw[0][2]),
    .data_o_gather_nw               (data_i_gather_nw[0][2]),
    .ready_i_gather_nw              (ready_o_gather_nw[0][2]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[0][2]),
    .data_i_merge_nw                (data_o_merge_nw[0][2]),
    .ready_o_merge_nw               (ready_i_merge_nw[0][2]),
    .valid_o_merge_nw               (valid_i_merge_nw[0][2]),
    .data_o_merge_nw                (data_i_merge_nw[0][2]),
    .ready_i_merge_nw               (ready_o_merge_nw[0][2]),

    .valid_i_cast_pe                (cast_valid_i_0_2),
    .data_i_cast_pe                 (cast_data_i_0_2),
    .ready_o_cast_pe                (cast_ready_o_0_2),
    .valid_o_cast_pe                (cast_valid_o_0_2),
    .data_o_cast_pe                 (cast_data_o_0_2),
    .ready_i_cast_pe                (cast_ready_i_0_2),

    .valid_i_merge_pe               (merge_valid_i_0_2),
    .data_i_merge_pe                (merge_data_i_0_2),
    .ready_o_merge_pe               (merge_ready_o_0_2),
    .valid_o_merge_pe               (merge_valid_o_0_2),
    .data_o_merge_pe                (merge_data_o_0_2),
    .ready_i_merge_pe               (merge_ready_i_0_2),

    .valid_i_gather_pe              (gather_valid_i_0_2),
    .data_i_gather_pe               (gather_data_i_0_2),
    .ready_o_gather_pe              (gather_ready_o_0_2),
    .valid_o_gather_pe              (gather_valid_o_0_2),
    .data_o_gather_pe               (gather_data_o_0_2),
    .ready_i_gather_pe              (gather_ready_i_0_2),

    .credit_upd                     (credit_upd[0][2])
);


network_interface #(
    .cast_out                       (cast_out_0_3),
    .gather_out                     (gather_out_0_3),
    .cast_sid                       (cast_sid_0_3),
    .gather_sid                     (gather_sid_0_3)
)ni_0_3(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[0][3]),
    .data_i_cast_nw                 (data_o_cast_nw[0][3]),
    .ready_o_cast_nw                (ready_i_cast_nw[0][3]),
    .valid_o_cast_nw                (valid_i_cast_nw[0][3]),
    .data_o_cast_nw                 (data_i_cast_nw[0][3]),
    .ready_i_cast_nw                (ready_o_cast_nw[0][3]),

    .valid_i_gather_nw              (valid_o_gather_nw[0][3]),
    .data_i_gather_nw               (data_o_gather_nw[0][3]),
    .ready_o_gather_nw              (ready_i_gather_nw[0][3]),
    .valid_o_gather_nw              (valid_i_gather_nw[0][3]),
    .data_o_gather_nw               (data_i_gather_nw[0][3]),
    .ready_i_gather_nw              (ready_o_gather_nw[0][3]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[0][3]),
    .data_i_merge_nw                (data_o_merge_nw[0][3]),
    .ready_o_merge_nw               (ready_i_merge_nw[0][3]),
    .valid_o_merge_nw               (valid_i_merge_nw[0][3]),
    .data_o_merge_nw                (data_i_merge_nw[0][3]),
    .ready_i_merge_nw               (ready_o_merge_nw[0][3]),

    .valid_i_cast_pe                (cast_valid_i_0_3),
    .data_i_cast_pe                 (cast_data_i_0_3),
    .ready_o_cast_pe                (cast_ready_o_0_3),
    .valid_o_cast_pe                (cast_valid_o_0_3),
    .data_o_cast_pe                 (cast_data_o_0_3),
    .ready_i_cast_pe                (cast_ready_i_0_3),

    .valid_i_merge_pe               (merge_valid_i_0_3),
    .data_i_merge_pe                (merge_data_i_0_3),
    .ready_o_merge_pe               (merge_ready_o_0_3),
    .valid_o_merge_pe               (merge_valid_o_0_3),
    .data_o_merge_pe                (merge_data_o_0_3),
    .ready_i_merge_pe               (merge_ready_i_0_3),

    .valid_i_gather_pe              (gather_valid_i_0_3),
    .data_i_gather_pe               (gather_data_i_0_3),
    .ready_o_gather_pe              (gather_ready_o_0_3),
    .valid_o_gather_pe              (gather_valid_o_0_3),
    .data_o_gather_pe               (gather_data_o_0_3),
    .ready_i_gather_pe              (gather_ready_i_0_3),

    .credit_upd                     (credit_upd[0][3])
);


network_interface #(
    .cast_out                       (cast_out_0_4),
    .gather_out                     (gather_out_0_4),
    .cast_sid                       (cast_sid_0_4),
    .gather_sid                     (gather_sid_0_4)
)ni_0_4(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[0][4]),
    .data_i_cast_nw                 (data_o_cast_nw[0][4]),
    .ready_o_cast_nw                (ready_i_cast_nw[0][4]),
    .valid_o_cast_nw                (valid_i_cast_nw[0][4]),
    .data_o_cast_nw                 (data_i_cast_nw[0][4]),
    .ready_i_cast_nw                (ready_o_cast_nw[0][4]),

    .valid_i_gather_nw              (valid_o_gather_nw[0][4]),
    .data_i_gather_nw               (data_o_gather_nw[0][4]),
    .ready_o_gather_nw              (ready_i_gather_nw[0][4]),
    .valid_o_gather_nw              (valid_i_gather_nw[0][4]),
    .data_o_gather_nw               (data_i_gather_nw[0][4]),
    .ready_i_gather_nw              (ready_o_gather_nw[0][4]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[0][4]),
    .data_i_merge_nw                (data_o_merge_nw[0][4]),
    .ready_o_merge_nw               (ready_i_merge_nw[0][4]),
    .valid_o_merge_nw               (valid_i_merge_nw[0][4]),
    .data_o_merge_nw                (data_i_merge_nw[0][4]),
    .ready_i_merge_nw               (ready_o_merge_nw[0][4]),

    .valid_i_cast_pe                (cast_valid_i_0_4),
    .data_i_cast_pe                 (cast_data_i_0_4),
    .ready_o_cast_pe                (cast_ready_o_0_4),
    .valid_o_cast_pe                (cast_valid_o_0_4),
    .data_o_cast_pe                 (cast_data_o_0_4),
    .ready_i_cast_pe                (cast_ready_i_0_4),

    .valid_i_merge_pe               (merge_valid_i_0_4),
    .data_i_merge_pe                (merge_data_i_0_4),
    .ready_o_merge_pe               (merge_ready_o_0_4),
    .valid_o_merge_pe               (merge_valid_o_0_4),
    .data_o_merge_pe                (merge_data_o_0_4),
    .ready_i_merge_pe               (merge_ready_i_0_4),

    .valid_i_gather_pe              (gather_valid_i_0_4),
    .data_i_gather_pe               (gather_data_i_0_4),
    .ready_o_gather_pe              (gather_ready_o_0_4),
    .valid_o_gather_pe              (gather_valid_o_0_4),
    .data_o_gather_pe               (gather_data_o_0_4),
    .ready_i_gather_pe              (gather_ready_i_0_4),

    .credit_upd                     (credit_upd[0][4])
);


network_interface #(
    .cast_out                       (cast_out_0_5),
    .gather_out                     (gather_out_0_5),
    .cast_sid                       (cast_sid_0_5),
    .gather_sid                     (gather_sid_0_5)
)ni_0_5(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[0][5]),
    .data_i_cast_nw                 (data_o_cast_nw[0][5]),
    .ready_o_cast_nw                (ready_i_cast_nw[0][5]),
    .valid_o_cast_nw                (valid_i_cast_nw[0][5]),
    .data_o_cast_nw                 (data_i_cast_nw[0][5]),
    .ready_i_cast_nw                (ready_o_cast_nw[0][5]),

    .valid_i_gather_nw              (valid_o_gather_nw[0][5]),
    .data_i_gather_nw               (data_o_gather_nw[0][5]),
    .ready_o_gather_nw              (ready_i_gather_nw[0][5]),
    .valid_o_gather_nw              (valid_i_gather_nw[0][5]),
    .data_o_gather_nw               (data_i_gather_nw[0][5]),
    .ready_i_gather_nw              (ready_o_gather_nw[0][5]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[0][5]),
    .data_i_merge_nw                (data_o_merge_nw[0][5]),
    .ready_o_merge_nw               (ready_i_merge_nw[0][5]),
    .valid_o_merge_nw               (valid_i_merge_nw[0][5]),
    .data_o_merge_nw                (data_i_merge_nw[0][5]),
    .ready_i_merge_nw               (ready_o_merge_nw[0][5]),

    .valid_i_cast_pe                (cast_valid_i_0_5),
    .data_i_cast_pe                 (cast_data_i_0_5),
    .ready_o_cast_pe                (cast_ready_o_0_5),
    .valid_o_cast_pe                (cast_valid_o_0_5),
    .data_o_cast_pe                 (cast_data_o_0_5),
    .ready_i_cast_pe                (cast_ready_i_0_5),

    .valid_i_merge_pe               (merge_valid_i_0_5),
    .data_i_merge_pe                (merge_data_i_0_5),
    .ready_o_merge_pe               (merge_ready_o_0_5),
    .valid_o_merge_pe               (merge_valid_o_0_5),
    .data_o_merge_pe                (merge_data_o_0_5),
    .ready_i_merge_pe               (merge_ready_i_0_5),

    .valid_i_gather_pe              (gather_valid_i_0_5),
    .data_i_gather_pe               (gather_data_i_0_5),
    .ready_o_gather_pe              (gather_ready_o_0_5),
    .valid_o_gather_pe              (gather_valid_o_0_5),
    .data_o_gather_pe               (gather_data_o_0_5),
    .ready_i_gather_pe              (gather_ready_i_0_5),

    .credit_upd                     (credit_upd[0][5])
);


network_interface #(
    .cast_out                       (cast_out_0_6),
    .gather_out                     (gather_out_0_6),
    .cast_sid                       (cast_sid_0_6),
    .gather_sid                     (gather_sid_0_6)
)ni_0_6(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[0][6]),
    .data_i_cast_nw                 (data_o_cast_nw[0][6]),
    .ready_o_cast_nw                (ready_i_cast_nw[0][6]),
    .valid_o_cast_nw                (valid_i_cast_nw[0][6]),
    .data_o_cast_nw                 (data_i_cast_nw[0][6]),
    .ready_i_cast_nw                (ready_o_cast_nw[0][6]),

    .valid_i_gather_nw              (valid_o_gather_nw[0][6]),
    .data_i_gather_nw               (data_o_gather_nw[0][6]),
    .ready_o_gather_nw              (ready_i_gather_nw[0][6]),
    .valid_o_gather_nw              (valid_i_gather_nw[0][6]),
    .data_o_gather_nw               (data_i_gather_nw[0][6]),
    .ready_i_gather_nw              (ready_o_gather_nw[0][6]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[0][6]),
    .data_i_merge_nw                (data_o_merge_nw[0][6]),
    .ready_o_merge_nw               (ready_i_merge_nw[0][6]),
    .valid_o_merge_nw               (valid_i_merge_nw[0][6]),
    .data_o_merge_nw                (data_i_merge_nw[0][6]),
    .ready_i_merge_nw               (ready_o_merge_nw[0][6]),

    .valid_i_cast_pe                (cast_valid_i_0_6),
    .data_i_cast_pe                 (cast_data_i_0_6),
    .ready_o_cast_pe                (cast_ready_o_0_6),
    .valid_o_cast_pe                (cast_valid_o_0_6),
    .data_o_cast_pe                 (cast_data_o_0_6),
    .ready_i_cast_pe                (cast_ready_i_0_6),

    .valid_i_merge_pe               (merge_valid_i_0_6),
    .data_i_merge_pe                (merge_data_i_0_6),
    .ready_o_merge_pe               (merge_ready_o_0_6),
    .valid_o_merge_pe               (merge_valid_o_0_6),
    .data_o_merge_pe                (merge_data_o_0_6),
    .ready_i_merge_pe               (merge_ready_i_0_6),

    .valid_i_gather_pe              (gather_valid_i_0_6),
    .data_i_gather_pe               (gather_data_i_0_6),
    .ready_o_gather_pe              (gather_ready_o_0_6),
    .valid_o_gather_pe              (gather_valid_o_0_6),
    .data_o_gather_pe               (gather_data_o_0_6),
    .ready_i_gather_pe              (gather_ready_i_0_6),

    .credit_upd                     (credit_upd[0][6])
);


network_interface #(
    .cast_out                       (cast_out_0_7),
    .gather_out                     (gather_out_0_7),
    .cast_sid                       (cast_sid_0_7),
    .gather_sid                     (gather_sid_0_7)
)ni_0_7(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[0][7]),
    .data_i_cast_nw                 (data_o_cast_nw[0][7]),
    .ready_o_cast_nw                (ready_i_cast_nw[0][7]),
    .valid_o_cast_nw                (valid_i_cast_nw[0][7]),
    .data_o_cast_nw                 (data_i_cast_nw[0][7]),
    .ready_i_cast_nw                (ready_o_cast_nw[0][7]),

    .valid_i_gather_nw              (valid_o_gather_nw[0][7]),
    .data_i_gather_nw               (data_o_gather_nw[0][7]),
    .ready_o_gather_nw              (ready_i_gather_nw[0][7]),
    .valid_o_gather_nw              (valid_i_gather_nw[0][7]),
    .data_o_gather_nw               (data_i_gather_nw[0][7]),
    .ready_i_gather_nw              (ready_o_gather_nw[0][7]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[0][7]),
    .data_i_merge_nw                (data_o_merge_nw[0][7]),
    .ready_o_merge_nw               (ready_i_merge_nw[0][7]),
    .valid_o_merge_nw               (valid_i_merge_nw[0][7]),
    .data_o_merge_nw                (data_i_merge_nw[0][7]),
    .ready_i_merge_nw               (ready_o_merge_nw[0][7]),

    .valid_i_cast_pe                (cast_valid_i_0_7),
    .data_i_cast_pe                 (cast_data_i_0_7),
    .ready_o_cast_pe                (cast_ready_o_0_7),
    .valid_o_cast_pe                (cast_valid_o_0_7),
    .data_o_cast_pe                 (cast_data_o_0_7),
    .ready_i_cast_pe                (cast_ready_i_0_7),

    .valid_i_merge_pe               (merge_valid_i_0_7),
    .data_i_merge_pe                (merge_data_i_0_7),
    .ready_o_merge_pe               (merge_ready_o_0_7),
    .valid_o_merge_pe               (merge_valid_o_0_7),
    .data_o_merge_pe                (merge_data_o_0_7),
    .ready_i_merge_pe               (merge_ready_i_0_7),

    .valid_i_gather_pe              (gather_valid_i_0_7),
    .data_i_gather_pe               (gather_data_i_0_7),
    .ready_o_gather_pe              (gather_ready_o_0_7),
    .valid_o_gather_pe              (gather_valid_o_0_7),
    .data_o_gather_pe               (gather_data_o_0_7),
    .ready_i_gather_pe              (gather_ready_i_0_7),

    .credit_upd                     (credit_upd[0][7])
);


network_interface #(
    .cast_out                       (cast_out_0_8),
    .gather_out                     (gather_out_0_8),
    .cast_sid                       (cast_sid_0_8),
    .gather_sid                     (gather_sid_0_8)
)ni_0_8(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[0][8]),
    .data_i_cast_nw                 (data_o_cast_nw[0][8]),
    .ready_o_cast_nw                (ready_i_cast_nw[0][8]),
    .valid_o_cast_nw                (valid_i_cast_nw[0][8]),
    .data_o_cast_nw                 (data_i_cast_nw[0][8]),
    .ready_i_cast_nw                (ready_o_cast_nw[0][8]),

    .valid_i_gather_nw              (valid_o_gather_nw[0][8]),
    .data_i_gather_nw               (data_o_gather_nw[0][8]),
    .ready_o_gather_nw              (ready_i_gather_nw[0][8]),
    .valid_o_gather_nw              (valid_i_gather_nw[0][8]),
    .data_o_gather_nw               (data_i_gather_nw[0][8]),
    .ready_i_gather_nw              (ready_o_gather_nw[0][8]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[0][8]),
    .data_i_merge_nw                (data_o_merge_nw[0][8]),
    .ready_o_merge_nw               (ready_i_merge_nw[0][8]),
    .valid_o_merge_nw               (valid_i_merge_nw[0][8]),
    .data_o_merge_nw                (data_i_merge_nw[0][8]),
    .ready_i_merge_nw               (ready_o_merge_nw[0][8]),

    .valid_i_cast_pe                (cast_valid_i_0_8),
    .data_i_cast_pe                 (cast_data_i_0_8),
    .ready_o_cast_pe                (cast_ready_o_0_8),
    .valid_o_cast_pe                (cast_valid_o_0_8),
    .data_o_cast_pe                 (cast_data_o_0_8),
    .ready_i_cast_pe                (cast_ready_i_0_8),

    .valid_i_merge_pe               (merge_valid_i_0_8),
    .data_i_merge_pe                (merge_data_i_0_8),
    .ready_o_merge_pe               (merge_ready_o_0_8),
    .valid_o_merge_pe               (merge_valid_o_0_8),
    .data_o_merge_pe                (merge_data_o_0_8),
    .ready_i_merge_pe               (merge_ready_i_0_8),

    .valid_i_gather_pe              (gather_valid_i_0_8),
    .data_i_gather_pe               (gather_data_i_0_8),
    .ready_o_gather_pe              (gather_ready_o_0_8),
    .valid_o_gather_pe              (gather_valid_o_0_8),
    .data_o_gather_pe               (gather_data_o_0_8),
    .ready_i_gather_pe              (gather_ready_i_0_8),

    .credit_upd                     (credit_upd[0][8])
);


network_interface #(
    .cast_out                       (cast_out_0_9),
    .gather_out                     (gather_out_0_9),
    .cast_sid                       (cast_sid_0_9),
    .gather_sid                     (gather_sid_0_9)
)ni_0_9(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[0][9]),
    .data_i_cast_nw                 (data_o_cast_nw[0][9]),
    .ready_o_cast_nw                (ready_i_cast_nw[0][9]),
    .valid_o_cast_nw                (valid_i_cast_nw[0][9]),
    .data_o_cast_nw                 (data_i_cast_nw[0][9]),
    .ready_i_cast_nw                (ready_o_cast_nw[0][9]),

    .valid_i_gather_nw              (valid_o_gather_nw[0][9]),
    .data_i_gather_nw               (data_o_gather_nw[0][9]),
    .ready_o_gather_nw              (ready_i_gather_nw[0][9]),
    .valid_o_gather_nw              (valid_i_gather_nw[0][9]),
    .data_o_gather_nw               (data_i_gather_nw[0][9]),
    .ready_i_gather_nw              (ready_o_gather_nw[0][9]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[0][9]),
    .data_i_merge_nw                (data_o_merge_nw[0][9]),
    .ready_o_merge_nw               (ready_i_merge_nw[0][9]),
    .valid_o_merge_nw               (valid_i_merge_nw[0][9]),
    .data_o_merge_nw                (data_i_merge_nw[0][9]),
    .ready_i_merge_nw               (ready_o_merge_nw[0][9]),

    .valid_i_cast_pe                (cast_valid_i_0_9),
    .data_i_cast_pe                 (cast_data_i_0_9),
    .ready_o_cast_pe                (cast_ready_o_0_9),
    .valid_o_cast_pe                (cast_valid_o_0_9),
    .data_o_cast_pe                 (cast_data_o_0_9),
    .ready_i_cast_pe                (cast_ready_i_0_9),

    .valid_i_merge_pe               (merge_valid_i_0_9),
    .data_i_merge_pe                (merge_data_i_0_9),
    .ready_o_merge_pe               (merge_ready_o_0_9),
    .valid_o_merge_pe               (merge_valid_o_0_9),
    .data_o_merge_pe                (merge_data_o_0_9),
    .ready_i_merge_pe               (merge_ready_i_0_9),

    .valid_i_gather_pe              (gather_valid_i_0_9),
    .data_i_gather_pe               (gather_data_i_0_9),
    .ready_o_gather_pe              (gather_ready_o_0_9),
    .valid_o_gather_pe              (gather_valid_o_0_9),
    .data_o_gather_pe               (gather_data_o_0_9),
    .ready_i_gather_pe              (gather_ready_i_0_9),

    .credit_upd                     (credit_upd[0][9])
);


network_interface #(
    .cast_out                       (cast_out_0_10),
    .gather_out                     (gather_out_0_10),
    .cast_sid                       (cast_sid_0_10),
    .gather_sid                     (gather_sid_0_10)
)ni_0_10(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[0][10]),
    .data_i_cast_nw                 (data_o_cast_nw[0][10]),
    .ready_o_cast_nw                (ready_i_cast_nw[0][10]),
    .valid_o_cast_nw                (valid_i_cast_nw[0][10]),
    .data_o_cast_nw                 (data_i_cast_nw[0][10]),
    .ready_i_cast_nw                (ready_o_cast_nw[0][10]),

    .valid_i_gather_nw              (valid_o_gather_nw[0][10]),
    .data_i_gather_nw               (data_o_gather_nw[0][10]),
    .ready_o_gather_nw              (ready_i_gather_nw[0][10]),
    .valid_o_gather_nw              (valid_i_gather_nw[0][10]),
    .data_o_gather_nw               (data_i_gather_nw[0][10]),
    .ready_i_gather_nw              (ready_o_gather_nw[0][10]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[0][10]),
    .data_i_merge_nw                (data_o_merge_nw[0][10]),
    .ready_o_merge_nw               (ready_i_merge_nw[0][10]),
    .valid_o_merge_nw               (valid_i_merge_nw[0][10]),
    .data_o_merge_nw                (data_i_merge_nw[0][10]),
    .ready_i_merge_nw               (ready_o_merge_nw[0][10]),

    .valid_i_cast_pe                (cast_valid_i_0_10),
    .data_i_cast_pe                 (cast_data_i_0_10),
    .ready_o_cast_pe                (cast_ready_o_0_10),
    .valid_o_cast_pe                (cast_valid_o_0_10),
    .data_o_cast_pe                 (cast_data_o_0_10),
    .ready_i_cast_pe                (cast_ready_i_0_10),

    .valid_i_merge_pe               (merge_valid_i_0_10),
    .data_i_merge_pe                (merge_data_i_0_10),
    .ready_o_merge_pe               (merge_ready_o_0_10),
    .valid_o_merge_pe               (merge_valid_o_0_10),
    .data_o_merge_pe                (merge_data_o_0_10),
    .ready_i_merge_pe               (merge_ready_i_0_10),

    .valid_i_gather_pe              (gather_valid_i_0_10),
    .data_i_gather_pe               (gather_data_i_0_10),
    .ready_o_gather_pe              (gather_ready_o_0_10),
    .valid_o_gather_pe              (gather_valid_o_0_10),
    .data_o_gather_pe               (gather_data_o_0_10),
    .ready_i_gather_pe              (gather_ready_i_0_10),

    .credit_upd                     (credit_upd[0][10])
);


network_interface #(
    .cast_out                       (cast_out_0_11),
    .gather_out                     (gather_out_0_11),
    .cast_sid                       (cast_sid_0_11),
    .gather_sid                     (gather_sid_0_11)
)ni_0_11(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[0][11]),
    .data_i_cast_nw                 (data_o_cast_nw[0][11]),
    .ready_o_cast_nw                (ready_i_cast_nw[0][11]),
    .valid_o_cast_nw                (valid_i_cast_nw[0][11]),
    .data_o_cast_nw                 (data_i_cast_nw[0][11]),
    .ready_i_cast_nw                (ready_o_cast_nw[0][11]),

    .valid_i_gather_nw              (valid_o_gather_nw[0][11]),
    .data_i_gather_nw               (data_o_gather_nw[0][11]),
    .ready_o_gather_nw              (ready_i_gather_nw[0][11]),
    .valid_o_gather_nw              (valid_i_gather_nw[0][11]),
    .data_o_gather_nw               (data_i_gather_nw[0][11]),
    .ready_i_gather_nw              (ready_o_gather_nw[0][11]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[0][11]),
    .data_i_merge_nw                (data_o_merge_nw[0][11]),
    .ready_o_merge_nw               (ready_i_merge_nw[0][11]),
    .valid_o_merge_nw               (valid_i_merge_nw[0][11]),
    .data_o_merge_nw                (data_i_merge_nw[0][11]),
    .ready_i_merge_nw               (ready_o_merge_nw[0][11]),

    .valid_i_cast_pe                (cast_valid_i_0_11),
    .data_i_cast_pe                 (cast_data_i_0_11),
    .ready_o_cast_pe                (cast_ready_o_0_11),
    .valid_o_cast_pe                (cast_valid_o_0_11),
    .data_o_cast_pe                 (cast_data_o_0_11),
    .ready_i_cast_pe                (cast_ready_i_0_11),

    .valid_i_merge_pe               (merge_valid_i_0_11),
    .data_i_merge_pe                (merge_data_i_0_11),
    .ready_o_merge_pe               (merge_ready_o_0_11),
    .valid_o_merge_pe               (merge_valid_o_0_11),
    .data_o_merge_pe                (merge_data_o_0_11),
    .ready_i_merge_pe               (merge_ready_i_0_11),

    .valid_i_gather_pe              (gather_valid_i_0_11),
    .data_i_gather_pe               (gather_data_i_0_11),
    .ready_o_gather_pe              (gather_ready_o_0_11),
    .valid_o_gather_pe              (gather_valid_o_0_11),
    .data_o_gather_pe               (gather_data_o_0_11),
    .ready_i_gather_pe              (gather_ready_i_0_11),

    .credit_upd                     (credit_upd[0][11])
);


network_interface #(
    .cast_out                       (cast_out_0_12),
    .gather_out                     (gather_out_0_12),
    .cast_sid                       (cast_sid_0_12),
    .gather_sid                     (gather_sid_0_12)
)ni_0_12(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[0][12]),
    .data_i_cast_nw                 (data_o_cast_nw[0][12]),
    .ready_o_cast_nw                (ready_i_cast_nw[0][12]),
    .valid_o_cast_nw                (valid_i_cast_nw[0][12]),
    .data_o_cast_nw                 (data_i_cast_nw[0][12]),
    .ready_i_cast_nw                (ready_o_cast_nw[0][12]),

    .valid_i_gather_nw              (valid_o_gather_nw[0][12]),
    .data_i_gather_nw               (data_o_gather_nw[0][12]),
    .ready_o_gather_nw              (ready_i_gather_nw[0][12]),
    .valid_o_gather_nw              (valid_i_gather_nw[0][12]),
    .data_o_gather_nw               (data_i_gather_nw[0][12]),
    .ready_i_gather_nw              (ready_o_gather_nw[0][12]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[0][12]),
    .data_i_merge_nw                (data_o_merge_nw[0][12]),
    .ready_o_merge_nw               (ready_i_merge_nw[0][12]),
    .valid_o_merge_nw               (valid_i_merge_nw[0][12]),
    .data_o_merge_nw                (data_i_merge_nw[0][12]),
    .ready_i_merge_nw               (ready_o_merge_nw[0][12]),

    .valid_i_cast_pe                (cast_valid_i_0_12),
    .data_i_cast_pe                 (cast_data_i_0_12),
    .ready_o_cast_pe                (cast_ready_o_0_12),
    .valid_o_cast_pe                (cast_valid_o_0_12),
    .data_o_cast_pe                 (cast_data_o_0_12),
    .ready_i_cast_pe                (cast_ready_i_0_12),

    .valid_i_merge_pe               (merge_valid_i_0_12),
    .data_i_merge_pe                (merge_data_i_0_12),
    .ready_o_merge_pe               (merge_ready_o_0_12),
    .valid_o_merge_pe               (merge_valid_o_0_12),
    .data_o_merge_pe                (merge_data_o_0_12),
    .ready_i_merge_pe               (merge_ready_i_0_12),

    .valid_i_gather_pe              (gather_valid_i_0_12),
    .data_i_gather_pe               (gather_data_i_0_12),
    .ready_o_gather_pe              (gather_ready_o_0_12),
    .valid_o_gather_pe              (gather_valid_o_0_12),
    .data_o_gather_pe               (gather_data_o_0_12),
    .ready_i_gather_pe              (gather_ready_i_0_12),

    .credit_upd                     (credit_upd[0][12])
);


network_interface #(
    .cast_out                       (cast_out_0_13),
    .gather_out                     (gather_out_0_13),
    .cast_sid                       (cast_sid_0_13),
    .gather_sid                     (gather_sid_0_13)
)ni_0_13(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[0][13]),
    .data_i_cast_nw                 (data_o_cast_nw[0][13]),
    .ready_o_cast_nw                (ready_i_cast_nw[0][13]),
    .valid_o_cast_nw                (valid_i_cast_nw[0][13]),
    .data_o_cast_nw                 (data_i_cast_nw[0][13]),
    .ready_i_cast_nw                (ready_o_cast_nw[0][13]),

    .valid_i_gather_nw              (valid_o_gather_nw[0][13]),
    .data_i_gather_nw               (data_o_gather_nw[0][13]),
    .ready_o_gather_nw              (ready_i_gather_nw[0][13]),
    .valid_o_gather_nw              (valid_i_gather_nw[0][13]),
    .data_o_gather_nw               (data_i_gather_nw[0][13]),
    .ready_i_gather_nw              (ready_o_gather_nw[0][13]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[0][13]),
    .data_i_merge_nw                (data_o_merge_nw[0][13]),
    .ready_o_merge_nw               (ready_i_merge_nw[0][13]),
    .valid_o_merge_nw               (valid_i_merge_nw[0][13]),
    .data_o_merge_nw                (data_i_merge_nw[0][13]),
    .ready_i_merge_nw               (ready_o_merge_nw[0][13]),

    .valid_i_cast_pe                (cast_valid_i_0_13),
    .data_i_cast_pe                 (cast_data_i_0_13),
    .ready_o_cast_pe                (cast_ready_o_0_13),
    .valid_o_cast_pe                (cast_valid_o_0_13),
    .data_o_cast_pe                 (cast_data_o_0_13),
    .ready_i_cast_pe                (cast_ready_i_0_13),

    .valid_i_merge_pe               (merge_valid_i_0_13),
    .data_i_merge_pe                (merge_data_i_0_13),
    .ready_o_merge_pe               (merge_ready_o_0_13),
    .valid_o_merge_pe               (merge_valid_o_0_13),
    .data_o_merge_pe                (merge_data_o_0_13),
    .ready_i_merge_pe               (merge_ready_i_0_13),

    .valid_i_gather_pe              (gather_valid_i_0_13),
    .data_i_gather_pe               (gather_data_i_0_13),
    .ready_o_gather_pe              (gather_ready_o_0_13),
    .valid_o_gather_pe              (gather_valid_o_0_13),
    .data_o_gather_pe               (gather_data_o_0_13),
    .ready_i_gather_pe              (gather_ready_i_0_13),

    .credit_upd                     (credit_upd[0][13])
);


network_interface #(
    .cast_out                       (cast_out_0_14),
    .gather_out                     (gather_out_0_14),
    .cast_sid                       (cast_sid_0_14),
    .gather_sid                     (gather_sid_0_14)
)ni_0_14(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[0][14]),
    .data_i_cast_nw                 (data_o_cast_nw[0][14]),
    .ready_o_cast_nw                (ready_i_cast_nw[0][14]),
    .valid_o_cast_nw                (valid_i_cast_nw[0][14]),
    .data_o_cast_nw                 (data_i_cast_nw[0][14]),
    .ready_i_cast_nw                (ready_o_cast_nw[0][14]),

    .valid_i_gather_nw              (valid_o_gather_nw[0][14]),
    .data_i_gather_nw               (data_o_gather_nw[0][14]),
    .ready_o_gather_nw              (ready_i_gather_nw[0][14]),
    .valid_o_gather_nw              (valid_i_gather_nw[0][14]),
    .data_o_gather_nw               (data_i_gather_nw[0][14]),
    .ready_i_gather_nw              (ready_o_gather_nw[0][14]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[0][14]),
    .data_i_merge_nw                (data_o_merge_nw[0][14]),
    .ready_o_merge_nw               (ready_i_merge_nw[0][14]),
    .valid_o_merge_nw               (valid_i_merge_nw[0][14]),
    .data_o_merge_nw                (data_i_merge_nw[0][14]),
    .ready_i_merge_nw               (ready_o_merge_nw[0][14]),

    .valid_i_cast_pe                (cast_valid_i_0_14),
    .data_i_cast_pe                 (cast_data_i_0_14),
    .ready_o_cast_pe                (cast_ready_o_0_14),
    .valid_o_cast_pe                (cast_valid_o_0_14),
    .data_o_cast_pe                 (cast_data_o_0_14),
    .ready_i_cast_pe                (cast_ready_i_0_14),

    .valid_i_merge_pe               (merge_valid_i_0_14),
    .data_i_merge_pe                (merge_data_i_0_14),
    .ready_o_merge_pe               (merge_ready_o_0_14),
    .valid_o_merge_pe               (merge_valid_o_0_14),
    .data_o_merge_pe                (merge_data_o_0_14),
    .ready_i_merge_pe               (merge_ready_i_0_14),

    .valid_i_gather_pe              (gather_valid_i_0_14),
    .data_i_gather_pe               (gather_data_i_0_14),
    .ready_o_gather_pe              (gather_ready_o_0_14),
    .valid_o_gather_pe              (gather_valid_o_0_14),
    .data_o_gather_pe               (gather_data_o_0_14),
    .ready_i_gather_pe              (gather_ready_i_0_14),

    .credit_upd                     (credit_upd[0][14])
);


network_interface #(
    .cast_out                       (cast_out_0_15),
    .gather_out                     (gather_out_0_15),
    .cast_sid                       (cast_sid_0_15),
    .gather_sid                     (gather_sid_0_15)
)ni_0_15(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[0][15]),
    .data_i_cast_nw                 (data_o_cast_nw[0][15]),
    .ready_o_cast_nw                (ready_i_cast_nw[0][15]),
    .valid_o_cast_nw                (valid_i_cast_nw[0][15]),
    .data_o_cast_nw                 (data_i_cast_nw[0][15]),
    .ready_i_cast_nw                (ready_o_cast_nw[0][15]),

    .valid_i_gather_nw              (valid_o_gather_nw[0][15]),
    .data_i_gather_nw               (data_o_gather_nw[0][15]),
    .ready_o_gather_nw              (ready_i_gather_nw[0][15]),
    .valid_o_gather_nw              (valid_i_gather_nw[0][15]),
    .data_o_gather_nw               (data_i_gather_nw[0][15]),
    .ready_i_gather_nw              (ready_o_gather_nw[0][15]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[0][15]),
    .data_i_merge_nw                (data_o_merge_nw[0][15]),
    .ready_o_merge_nw               (ready_i_merge_nw[0][15]),
    .valid_o_merge_nw               (valid_i_merge_nw[0][15]),
    .data_o_merge_nw                (data_i_merge_nw[0][15]),
    .ready_i_merge_nw               (ready_o_merge_nw[0][15]),

    .valid_i_cast_pe                (cast_valid_i_0_15),
    .data_i_cast_pe                 (cast_data_i_0_15),
    .ready_o_cast_pe                (cast_ready_o_0_15),
    .valid_o_cast_pe                (cast_valid_o_0_15),
    .data_o_cast_pe                 (cast_data_o_0_15),
    .ready_i_cast_pe                (cast_ready_i_0_15),

    .valid_i_merge_pe               (merge_valid_i_0_15),
    .data_i_merge_pe                (merge_data_i_0_15),
    .ready_o_merge_pe               (merge_ready_o_0_15),
    .valid_o_merge_pe               (merge_valid_o_0_15),
    .data_o_merge_pe                (merge_data_o_0_15),
    .ready_i_merge_pe               (merge_ready_i_0_15),

    .valid_i_gather_pe              (gather_valid_i_0_15),
    .data_i_gather_pe               (gather_data_i_0_15),
    .ready_o_gather_pe              (gather_ready_o_0_15),
    .valid_o_gather_pe              (gather_valid_o_0_15),
    .data_o_gather_pe               (gather_data_o_0_15),
    .ready_i_gather_pe              (gather_ready_i_0_15),

    .credit_upd                     (credit_upd[0][15])
);


network_interface #(
    .cast_out                       (cast_out_0_16),
    .gather_out                     (gather_out_0_16),
    .cast_sid                       (cast_sid_0_16),
    .gather_sid                     (gather_sid_0_16)
)ni_0_16(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[0][16]),
    .data_i_cast_nw                 (data_o_cast_nw[0][16]),
    .ready_o_cast_nw                (ready_i_cast_nw[0][16]),
    .valid_o_cast_nw                (valid_i_cast_nw[0][16]),
    .data_o_cast_nw                 (data_i_cast_nw[0][16]),
    .ready_i_cast_nw                (ready_o_cast_nw[0][16]),

    .valid_i_gather_nw              (valid_o_gather_nw[0][16]),
    .data_i_gather_nw               (data_o_gather_nw[0][16]),
    .ready_o_gather_nw              (ready_i_gather_nw[0][16]),
    .valid_o_gather_nw              (valid_i_gather_nw[0][16]),
    .data_o_gather_nw               (data_i_gather_nw[0][16]),
    .ready_i_gather_nw              (ready_o_gather_nw[0][16]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[0][16]),
    .data_i_merge_nw                (data_o_merge_nw[0][16]),
    .ready_o_merge_nw               (ready_i_merge_nw[0][16]),
    .valid_o_merge_nw               (valid_i_merge_nw[0][16]),
    .data_o_merge_nw                (data_i_merge_nw[0][16]),
    .ready_i_merge_nw               (ready_o_merge_nw[0][16]),

    .valid_i_cast_pe                (cast_valid_i_0_16),
    .data_i_cast_pe                 (cast_data_i_0_16),
    .ready_o_cast_pe                (cast_ready_o_0_16),
    .valid_o_cast_pe                (cast_valid_o_0_16),
    .data_o_cast_pe                 (cast_data_o_0_16),
    .ready_i_cast_pe                (cast_ready_i_0_16),

    .valid_i_merge_pe               (merge_valid_i_0_16),
    .data_i_merge_pe                (merge_data_i_0_16),
    .ready_o_merge_pe               (merge_ready_o_0_16),
    .valid_o_merge_pe               (merge_valid_o_0_16),
    .data_o_merge_pe                (merge_data_o_0_16),
    .ready_i_merge_pe               (merge_ready_i_0_16),

    .valid_i_gather_pe              (gather_valid_i_0_16),
    .data_i_gather_pe               (gather_data_i_0_16),
    .ready_o_gather_pe              (gather_ready_o_0_16),
    .valid_o_gather_pe              (gather_valid_o_0_16),
    .data_o_gather_pe               (gather_data_o_0_16),
    .ready_i_gather_pe              (gather_ready_i_0_16),

    .credit_upd                     (credit_upd[0][16])
);


network_interface #(
    .cast_out                       (cast_out_0_17),
    .gather_out                     (gather_out_0_17),
    .cast_sid                       (cast_sid_0_17),
    .gather_sid                     (gather_sid_0_17)
)ni_0_17(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[0][17]),
    .data_i_cast_nw                 (data_o_cast_nw[0][17]),
    .ready_o_cast_nw                (ready_i_cast_nw[0][17]),
    .valid_o_cast_nw                (valid_i_cast_nw[0][17]),
    .data_o_cast_nw                 (data_i_cast_nw[0][17]),
    .ready_i_cast_nw                (ready_o_cast_nw[0][17]),

    .valid_i_gather_nw              (valid_o_gather_nw[0][17]),
    .data_i_gather_nw               (data_o_gather_nw[0][17]),
    .ready_o_gather_nw              (ready_i_gather_nw[0][17]),
    .valid_o_gather_nw              (valid_i_gather_nw[0][17]),
    .data_o_gather_nw               (data_i_gather_nw[0][17]),
    .ready_i_gather_nw              (ready_o_gather_nw[0][17]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[0][17]),
    .data_i_merge_nw                (data_o_merge_nw[0][17]),
    .ready_o_merge_nw               (ready_i_merge_nw[0][17]),
    .valid_o_merge_nw               (valid_i_merge_nw[0][17]),
    .data_o_merge_nw                (data_i_merge_nw[0][17]),
    .ready_i_merge_nw               (ready_o_merge_nw[0][17]),

    .valid_i_cast_pe                (cast_valid_i_0_17),
    .data_i_cast_pe                 (cast_data_i_0_17),
    .ready_o_cast_pe                (cast_ready_o_0_17),
    .valid_o_cast_pe                (cast_valid_o_0_17),
    .data_o_cast_pe                 (cast_data_o_0_17),
    .ready_i_cast_pe                (cast_ready_i_0_17),

    .valid_i_merge_pe               (merge_valid_i_0_17),
    .data_i_merge_pe                (merge_data_i_0_17),
    .ready_o_merge_pe               (merge_ready_o_0_17),
    .valid_o_merge_pe               (merge_valid_o_0_17),
    .data_o_merge_pe                (merge_data_o_0_17),
    .ready_i_merge_pe               (merge_ready_i_0_17),

    .valid_i_gather_pe              (gather_valid_i_0_17),
    .data_i_gather_pe               (gather_data_i_0_17),
    .ready_o_gather_pe              (gather_ready_o_0_17),
    .valid_o_gather_pe              (gather_valid_o_0_17),
    .data_o_gather_pe               (gather_data_o_0_17),
    .ready_i_gather_pe              (gather_ready_i_0_17),

    .credit_upd                     (credit_upd[0][17])
);


network_interface #(
    .cast_out                       (cast_out_0_18),
    .gather_out                     (gather_out_0_18),
    .cast_sid                       (cast_sid_0_18),
    .gather_sid                     (gather_sid_0_18)
)ni_0_18(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[0][18]),
    .data_i_cast_nw                 (data_o_cast_nw[0][18]),
    .ready_o_cast_nw                (ready_i_cast_nw[0][18]),
    .valid_o_cast_nw                (valid_i_cast_nw[0][18]),
    .data_o_cast_nw                 (data_i_cast_nw[0][18]),
    .ready_i_cast_nw                (ready_o_cast_nw[0][18]),

    .valid_i_gather_nw              (valid_o_gather_nw[0][18]),
    .data_i_gather_nw               (data_o_gather_nw[0][18]),
    .ready_o_gather_nw              (ready_i_gather_nw[0][18]),
    .valid_o_gather_nw              (valid_i_gather_nw[0][18]),
    .data_o_gather_nw               (data_i_gather_nw[0][18]),
    .ready_i_gather_nw              (ready_o_gather_nw[0][18]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[0][18]),
    .data_i_merge_nw                (data_o_merge_nw[0][18]),
    .ready_o_merge_nw               (ready_i_merge_nw[0][18]),
    .valid_o_merge_nw               (valid_i_merge_nw[0][18]),
    .data_o_merge_nw                (data_i_merge_nw[0][18]),
    .ready_i_merge_nw               (ready_o_merge_nw[0][18]),

    .valid_i_cast_pe                (cast_valid_i_0_18),
    .data_i_cast_pe                 (cast_data_i_0_18),
    .ready_o_cast_pe                (cast_ready_o_0_18),
    .valid_o_cast_pe                (cast_valid_o_0_18),
    .data_o_cast_pe                 (cast_data_o_0_18),
    .ready_i_cast_pe                (cast_ready_i_0_18),

    .valid_i_merge_pe               (merge_valid_i_0_18),
    .data_i_merge_pe                (merge_data_i_0_18),
    .ready_o_merge_pe               (merge_ready_o_0_18),
    .valid_o_merge_pe               (merge_valid_o_0_18),
    .data_o_merge_pe                (merge_data_o_0_18),
    .ready_i_merge_pe               (merge_ready_i_0_18),

    .valid_i_gather_pe              (gather_valid_i_0_18),
    .data_i_gather_pe               (gather_data_i_0_18),
    .ready_o_gather_pe              (gather_ready_o_0_18),
    .valid_o_gather_pe              (gather_valid_o_0_18),
    .data_o_gather_pe               (gather_data_o_0_18),
    .ready_i_gather_pe              (gather_ready_i_0_18),

    .credit_upd                     (credit_upd[0][18])
);


network_interface #(
    .cast_out                       (cast_out_0_19),
    .gather_out                     (gather_out_0_19),
    .cast_sid                       (cast_sid_0_19),
    .gather_sid                     (gather_sid_0_19)
)ni_0_19(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[0][19]),
    .data_i_cast_nw                 (data_o_cast_nw[0][19]),
    .ready_o_cast_nw                (ready_i_cast_nw[0][19]),
    .valid_o_cast_nw                (valid_i_cast_nw[0][19]),
    .data_o_cast_nw                 (data_i_cast_nw[0][19]),
    .ready_i_cast_nw                (ready_o_cast_nw[0][19]),

    .valid_i_gather_nw              (valid_o_gather_nw[0][19]),
    .data_i_gather_nw               (data_o_gather_nw[0][19]),
    .ready_o_gather_nw              (ready_i_gather_nw[0][19]),
    .valid_o_gather_nw              (valid_i_gather_nw[0][19]),
    .data_o_gather_nw               (data_i_gather_nw[0][19]),
    .ready_i_gather_nw              (ready_o_gather_nw[0][19]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[0][19]),
    .data_i_merge_nw                (data_o_merge_nw[0][19]),
    .ready_o_merge_nw               (ready_i_merge_nw[0][19]),
    .valid_o_merge_nw               (valid_i_merge_nw[0][19]),
    .data_o_merge_nw                (data_i_merge_nw[0][19]),
    .ready_i_merge_nw               (ready_o_merge_nw[0][19]),

    .valid_i_cast_pe                (cast_valid_i_0_19),
    .data_i_cast_pe                 (cast_data_i_0_19),
    .ready_o_cast_pe                (cast_ready_o_0_19),
    .valid_o_cast_pe                (cast_valid_o_0_19),
    .data_o_cast_pe                 (cast_data_o_0_19),
    .ready_i_cast_pe                (cast_ready_i_0_19),

    .valid_i_merge_pe               (merge_valid_i_0_19),
    .data_i_merge_pe                (merge_data_i_0_19),
    .ready_o_merge_pe               (merge_ready_o_0_19),
    .valid_o_merge_pe               (merge_valid_o_0_19),
    .data_o_merge_pe                (merge_data_o_0_19),
    .ready_i_merge_pe               (merge_ready_i_0_19),

    .valid_i_gather_pe              (gather_valid_i_0_19),
    .data_i_gather_pe               (gather_data_i_0_19),
    .ready_o_gather_pe              (gather_ready_o_0_19),
    .valid_o_gather_pe              (gather_valid_o_0_19),
    .data_o_gather_pe               (gather_data_o_0_19),
    .ready_i_gather_pe              (gather_ready_i_0_19),

    .credit_upd                     (credit_upd[0][19])
);


network_interface #(
    .cast_out                       (cast_out_0_20),
    .gather_out                     (gather_out_0_20),
    .cast_sid                       (cast_sid_0_20),
    .gather_sid                     (gather_sid_0_20)
)ni_0_20(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[0][20]),
    .data_i_cast_nw                 (data_o_cast_nw[0][20]),
    .ready_o_cast_nw                (ready_i_cast_nw[0][20]),
    .valid_o_cast_nw                (valid_i_cast_nw[0][20]),
    .data_o_cast_nw                 (data_i_cast_nw[0][20]),
    .ready_i_cast_nw                (ready_o_cast_nw[0][20]),

    .valid_i_gather_nw              (valid_o_gather_nw[0][20]),
    .data_i_gather_nw               (data_o_gather_nw[0][20]),
    .ready_o_gather_nw              (ready_i_gather_nw[0][20]),
    .valid_o_gather_nw              (valid_i_gather_nw[0][20]),
    .data_o_gather_nw               (data_i_gather_nw[0][20]),
    .ready_i_gather_nw              (ready_o_gather_nw[0][20]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[0][20]),
    .data_i_merge_nw                (data_o_merge_nw[0][20]),
    .ready_o_merge_nw               (ready_i_merge_nw[0][20]),
    .valid_o_merge_nw               (valid_i_merge_nw[0][20]),
    .data_o_merge_nw                (data_i_merge_nw[0][20]),
    .ready_i_merge_nw               (ready_o_merge_nw[0][20]),

    .valid_i_cast_pe                (cast_valid_i_0_20),
    .data_i_cast_pe                 (cast_data_i_0_20),
    .ready_o_cast_pe                (cast_ready_o_0_20),
    .valid_o_cast_pe                (cast_valid_o_0_20),
    .data_o_cast_pe                 (cast_data_o_0_20),
    .ready_i_cast_pe                (cast_ready_i_0_20),

    .valid_i_merge_pe               (merge_valid_i_0_20),
    .data_i_merge_pe                (merge_data_i_0_20),
    .ready_o_merge_pe               (merge_ready_o_0_20),
    .valid_o_merge_pe               (merge_valid_o_0_20),
    .data_o_merge_pe                (merge_data_o_0_20),
    .ready_i_merge_pe               (merge_ready_i_0_20),

    .valid_i_gather_pe              (gather_valid_i_0_20),
    .data_i_gather_pe               (gather_data_i_0_20),
    .ready_o_gather_pe              (gather_ready_o_0_20),
    .valid_o_gather_pe              (gather_valid_o_0_20),
    .data_o_gather_pe               (gather_data_o_0_20),
    .ready_i_gather_pe              (gather_ready_i_0_20),

    .credit_upd                     (credit_upd[0][20])
);


network_interface #(
    .cast_out                       (cast_out_0_21),
    .gather_out                     (gather_out_0_21),
    .cast_sid                       (cast_sid_0_21),
    .gather_sid                     (gather_sid_0_21)
)ni_0_21(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[0][21]),
    .data_i_cast_nw                 (data_o_cast_nw[0][21]),
    .ready_o_cast_nw                (ready_i_cast_nw[0][21]),
    .valid_o_cast_nw                (valid_i_cast_nw[0][21]),
    .data_o_cast_nw                 (data_i_cast_nw[0][21]),
    .ready_i_cast_nw                (ready_o_cast_nw[0][21]),

    .valid_i_gather_nw              (valid_o_gather_nw[0][21]),
    .data_i_gather_nw               (data_o_gather_nw[0][21]),
    .ready_o_gather_nw              (ready_i_gather_nw[0][21]),
    .valid_o_gather_nw              (valid_i_gather_nw[0][21]),
    .data_o_gather_nw               (data_i_gather_nw[0][21]),
    .ready_i_gather_nw              (ready_o_gather_nw[0][21]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[0][21]),
    .data_i_merge_nw                (data_o_merge_nw[0][21]),
    .ready_o_merge_nw               (ready_i_merge_nw[0][21]),
    .valid_o_merge_nw               (valid_i_merge_nw[0][21]),
    .data_o_merge_nw                (data_i_merge_nw[0][21]),
    .ready_i_merge_nw               (ready_o_merge_nw[0][21]),

    .valid_i_cast_pe                (cast_valid_i_0_21),
    .data_i_cast_pe                 (cast_data_i_0_21),
    .ready_o_cast_pe                (cast_ready_o_0_21),
    .valid_o_cast_pe                (cast_valid_o_0_21),
    .data_o_cast_pe                 (cast_data_o_0_21),
    .ready_i_cast_pe                (cast_ready_i_0_21),

    .valid_i_merge_pe               (merge_valid_i_0_21),
    .data_i_merge_pe                (merge_data_i_0_21),
    .ready_o_merge_pe               (merge_ready_o_0_21),
    .valid_o_merge_pe               (merge_valid_o_0_21),
    .data_o_merge_pe                (merge_data_o_0_21),
    .ready_i_merge_pe               (merge_ready_i_0_21),

    .valid_i_gather_pe              (gather_valid_i_0_21),
    .data_i_gather_pe               (gather_data_i_0_21),
    .ready_o_gather_pe              (gather_ready_o_0_21),
    .valid_o_gather_pe              (gather_valid_o_0_21),
    .data_o_gather_pe               (gather_data_o_0_21),
    .ready_i_gather_pe              (gather_ready_i_0_21),

    .credit_upd                     (credit_upd[0][21])
);


network_interface #(
    .cast_out                       (cast_out_0_22),
    .gather_out                     (gather_out_0_22),
    .cast_sid                       (cast_sid_0_22),
    .gather_sid                     (gather_sid_0_22)
)ni_0_22(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[0][22]),
    .data_i_cast_nw                 (data_o_cast_nw[0][22]),
    .ready_o_cast_nw                (ready_i_cast_nw[0][22]),
    .valid_o_cast_nw                (valid_i_cast_nw[0][22]),
    .data_o_cast_nw                 (data_i_cast_nw[0][22]),
    .ready_i_cast_nw                (ready_o_cast_nw[0][22]),

    .valid_i_gather_nw              (valid_o_gather_nw[0][22]),
    .data_i_gather_nw               (data_o_gather_nw[0][22]),
    .ready_o_gather_nw              (ready_i_gather_nw[0][22]),
    .valid_o_gather_nw              (valid_i_gather_nw[0][22]),
    .data_o_gather_nw               (data_i_gather_nw[0][22]),
    .ready_i_gather_nw              (ready_o_gather_nw[0][22]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[0][22]),
    .data_i_merge_nw                (data_o_merge_nw[0][22]),
    .ready_o_merge_nw               (ready_i_merge_nw[0][22]),
    .valid_o_merge_nw               (valid_i_merge_nw[0][22]),
    .data_o_merge_nw                (data_i_merge_nw[0][22]),
    .ready_i_merge_nw               (ready_o_merge_nw[0][22]),

    .valid_i_cast_pe                (cast_valid_i_0_22),
    .data_i_cast_pe                 (cast_data_i_0_22),
    .ready_o_cast_pe                (cast_ready_o_0_22),
    .valid_o_cast_pe                (cast_valid_o_0_22),
    .data_o_cast_pe                 (cast_data_o_0_22),
    .ready_i_cast_pe                (cast_ready_i_0_22),

    .valid_i_merge_pe               (merge_valid_i_0_22),
    .data_i_merge_pe                (merge_data_i_0_22),
    .ready_o_merge_pe               (merge_ready_o_0_22),
    .valid_o_merge_pe               (merge_valid_o_0_22),
    .data_o_merge_pe                (merge_data_o_0_22),
    .ready_i_merge_pe               (merge_ready_i_0_22),

    .valid_i_gather_pe              (gather_valid_i_0_22),
    .data_i_gather_pe               (gather_data_i_0_22),
    .ready_o_gather_pe              (gather_ready_o_0_22),
    .valid_o_gather_pe              (gather_valid_o_0_22),
    .data_o_gather_pe               (gather_data_o_0_22),
    .ready_i_gather_pe              (gather_ready_i_0_22),

    .credit_upd                     (credit_upd[0][22])
);


network_interface #(
    .cast_out                       (cast_out_0_23),
    .gather_out                     (gather_out_0_23),
    .cast_sid                       (cast_sid_0_23),
    .gather_sid                     (gather_sid_0_23)
)ni_0_23(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[0][23]),
    .data_i_cast_nw                 (data_o_cast_nw[0][23]),
    .ready_o_cast_nw                (ready_i_cast_nw[0][23]),
    .valid_o_cast_nw                (valid_i_cast_nw[0][23]),
    .data_o_cast_nw                 (data_i_cast_nw[0][23]),
    .ready_i_cast_nw                (ready_o_cast_nw[0][23]),

    .valid_i_gather_nw              (valid_o_gather_nw[0][23]),
    .data_i_gather_nw               (data_o_gather_nw[0][23]),
    .ready_o_gather_nw              (ready_i_gather_nw[0][23]),
    .valid_o_gather_nw              (valid_i_gather_nw[0][23]),
    .data_o_gather_nw               (data_i_gather_nw[0][23]),
    .ready_i_gather_nw              (ready_o_gather_nw[0][23]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[0][23]),
    .data_i_merge_nw                (data_o_merge_nw[0][23]),
    .ready_o_merge_nw               (ready_i_merge_nw[0][23]),
    .valid_o_merge_nw               (valid_i_merge_nw[0][23]),
    .data_o_merge_nw                (data_i_merge_nw[0][23]),
    .ready_i_merge_nw               (ready_o_merge_nw[0][23]),

    .valid_i_cast_pe                (cast_valid_i_0_23),
    .data_i_cast_pe                 (cast_data_i_0_23),
    .ready_o_cast_pe                (cast_ready_o_0_23),
    .valid_o_cast_pe                (cast_valid_o_0_23),
    .data_o_cast_pe                 (cast_data_o_0_23),
    .ready_i_cast_pe                (cast_ready_i_0_23),

    .valid_i_merge_pe               (merge_valid_i_0_23),
    .data_i_merge_pe                (merge_data_i_0_23),
    .ready_o_merge_pe               (merge_ready_o_0_23),
    .valid_o_merge_pe               (merge_valid_o_0_23),
    .data_o_merge_pe                (merge_data_o_0_23),
    .ready_i_merge_pe               (merge_ready_i_0_23),

    .valid_i_gather_pe              (gather_valid_i_0_23),
    .data_i_gather_pe               (gather_data_i_0_23),
    .ready_o_gather_pe              (gather_ready_o_0_23),
    .valid_o_gather_pe              (gather_valid_o_0_23),
    .data_o_gather_pe               (gather_data_o_0_23),
    .ready_i_gather_pe              (gather_ready_i_0_23),

    .credit_upd                     (credit_upd[0][23])
);


network_interface #(
    .cast_out                       (cast_out_0_24),
    .gather_out                     (gather_out_0_24),
    .cast_sid                       (cast_sid_0_24),
    .gather_sid                     (gather_sid_0_24)
)ni_0_24(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[0][24]),
    .data_i_cast_nw                 (data_o_cast_nw[0][24]),
    .ready_o_cast_nw                (ready_i_cast_nw[0][24]),
    .valid_o_cast_nw                (valid_i_cast_nw[0][24]),
    .data_o_cast_nw                 (data_i_cast_nw[0][24]),
    .ready_i_cast_nw                (ready_o_cast_nw[0][24]),

    .valid_i_gather_nw              (valid_o_gather_nw[0][24]),
    .data_i_gather_nw               (data_o_gather_nw[0][24]),
    .ready_o_gather_nw              (ready_i_gather_nw[0][24]),
    .valid_o_gather_nw              (valid_i_gather_nw[0][24]),
    .data_o_gather_nw               (data_i_gather_nw[0][24]),
    .ready_i_gather_nw              (ready_o_gather_nw[0][24]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[0][24]),
    .data_i_merge_nw                (data_o_merge_nw[0][24]),
    .ready_o_merge_nw               (ready_i_merge_nw[0][24]),
    .valid_o_merge_nw               (valid_i_merge_nw[0][24]),
    .data_o_merge_nw                (data_i_merge_nw[0][24]),
    .ready_i_merge_nw               (ready_o_merge_nw[0][24]),

    .valid_i_cast_pe                (cast_valid_i_0_24),
    .data_i_cast_pe                 (cast_data_i_0_24),
    .ready_o_cast_pe                (cast_ready_o_0_24),
    .valid_o_cast_pe                (cast_valid_o_0_24),
    .data_o_cast_pe                 (cast_data_o_0_24),
    .ready_i_cast_pe                (cast_ready_i_0_24),

    .valid_i_merge_pe               (merge_valid_i_0_24),
    .data_i_merge_pe                (merge_data_i_0_24),
    .ready_o_merge_pe               (merge_ready_o_0_24),
    .valid_o_merge_pe               (merge_valid_o_0_24),
    .data_o_merge_pe                (merge_data_o_0_24),
    .ready_i_merge_pe               (merge_ready_i_0_24),

    .valid_i_gather_pe              (gather_valid_i_0_24),
    .data_i_gather_pe               (gather_data_i_0_24),
    .ready_o_gather_pe              (gather_ready_o_0_24),
    .valid_o_gather_pe              (gather_valid_o_0_24),
    .data_o_gather_pe               (gather_data_o_0_24),
    .ready_i_gather_pe              (gather_ready_i_0_24),

    .credit_upd                     (credit_upd[0][24])
);


network_interface #(
    .cast_out                       (cast_out_1_0),
    .gather_out                     (gather_out_1_0),
    .cast_sid                       (cast_sid_1_0),
    .gather_sid                     (gather_sid_1_0)
)ni_1_0(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[1][0]),
    .data_i_cast_nw                 (data_o_cast_nw[1][0]),
    .ready_o_cast_nw                (ready_i_cast_nw[1][0]),
    .valid_o_cast_nw                (valid_i_cast_nw[1][0]),
    .data_o_cast_nw                 (data_i_cast_nw[1][0]),
    .ready_i_cast_nw                (ready_o_cast_nw[1][0]),

    .valid_i_gather_nw              (valid_o_gather_nw[1][0]),
    .data_i_gather_nw               (data_o_gather_nw[1][0]),
    .ready_o_gather_nw              (ready_i_gather_nw[1][0]),
    .valid_o_gather_nw              (valid_i_gather_nw[1][0]),
    .data_o_gather_nw               (data_i_gather_nw[1][0]),
    .ready_i_gather_nw              (ready_o_gather_nw[1][0]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[1][0]),
    .data_i_merge_nw                (data_o_merge_nw[1][0]),
    .ready_o_merge_nw               (ready_i_merge_nw[1][0]),
    .valid_o_merge_nw               (valid_i_merge_nw[1][0]),
    .data_o_merge_nw                (data_i_merge_nw[1][0]),
    .ready_i_merge_nw               (ready_o_merge_nw[1][0]),

    .valid_i_cast_pe                (cast_valid_i_1_0),
    .data_i_cast_pe                 (cast_data_i_1_0),
    .ready_o_cast_pe                (cast_ready_o_1_0),
    .valid_o_cast_pe                (cast_valid_o_1_0),
    .data_o_cast_pe                 (cast_data_o_1_0),
    .ready_i_cast_pe                (cast_ready_i_1_0),

    .valid_i_merge_pe               (merge_valid_i_1_0),
    .data_i_merge_pe                (merge_data_i_1_0),
    .ready_o_merge_pe               (merge_ready_o_1_0),
    .valid_o_merge_pe               (merge_valid_o_1_0),
    .data_o_merge_pe                (merge_data_o_1_0),
    .ready_i_merge_pe               (merge_ready_i_1_0),

    .valid_i_gather_pe              (gather_valid_i_1_0),
    .data_i_gather_pe               (gather_data_i_1_0),
    .ready_o_gather_pe              (gather_ready_o_1_0),
    .valid_o_gather_pe              (gather_valid_o_1_0),
    .data_o_gather_pe               (gather_data_o_1_0),
    .ready_i_gather_pe              (gather_ready_i_1_0),

    .credit_upd                     (credit_upd[1][0])
);


network_interface #(
    .cast_out                       (cast_out_1_1),
    .gather_out                     (gather_out_1_1),
    .cast_sid                       (cast_sid_1_1),
    .gather_sid                     (gather_sid_1_1)
)ni_1_1(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[1][1]),
    .data_i_cast_nw                 (data_o_cast_nw[1][1]),
    .ready_o_cast_nw                (ready_i_cast_nw[1][1]),
    .valid_o_cast_nw                (valid_i_cast_nw[1][1]),
    .data_o_cast_nw                 (data_i_cast_nw[1][1]),
    .ready_i_cast_nw                (ready_o_cast_nw[1][1]),

    .valid_i_gather_nw              (valid_o_gather_nw[1][1]),
    .data_i_gather_nw               (data_o_gather_nw[1][1]),
    .ready_o_gather_nw              (ready_i_gather_nw[1][1]),
    .valid_o_gather_nw              (valid_i_gather_nw[1][1]),
    .data_o_gather_nw               (data_i_gather_nw[1][1]),
    .ready_i_gather_nw              (ready_o_gather_nw[1][1]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[1][1]),
    .data_i_merge_nw                (data_o_merge_nw[1][1]),
    .ready_o_merge_nw               (ready_i_merge_nw[1][1]),
    .valid_o_merge_nw               (valid_i_merge_nw[1][1]),
    .data_o_merge_nw                (data_i_merge_nw[1][1]),
    .ready_i_merge_nw               (ready_o_merge_nw[1][1]),

    .valid_i_cast_pe                (cast_valid_i_1_1),
    .data_i_cast_pe                 (cast_data_i_1_1),
    .ready_o_cast_pe                (cast_ready_o_1_1),
    .valid_o_cast_pe                (cast_valid_o_1_1),
    .data_o_cast_pe                 (cast_data_o_1_1),
    .ready_i_cast_pe                (cast_ready_i_1_1),

    .valid_i_merge_pe               (merge_valid_i_1_1),
    .data_i_merge_pe                (merge_data_i_1_1),
    .ready_o_merge_pe               (merge_ready_o_1_1),
    .valid_o_merge_pe               (merge_valid_o_1_1),
    .data_o_merge_pe                (merge_data_o_1_1),
    .ready_i_merge_pe               (merge_ready_i_1_1),

    .valid_i_gather_pe              (gather_valid_i_1_1),
    .data_i_gather_pe               (gather_data_i_1_1),
    .ready_o_gather_pe              (gather_ready_o_1_1),
    .valid_o_gather_pe              (gather_valid_o_1_1),
    .data_o_gather_pe               (gather_data_o_1_1),
    .ready_i_gather_pe              (gather_ready_i_1_1),

    .credit_upd                     (credit_upd[1][1])
);


network_interface #(
    .cast_out                       (cast_out_1_2),
    .gather_out                     (gather_out_1_2),
    .cast_sid                       (cast_sid_1_2),
    .gather_sid                     (gather_sid_1_2)
)ni_1_2(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[1][2]),
    .data_i_cast_nw                 (data_o_cast_nw[1][2]),
    .ready_o_cast_nw                (ready_i_cast_nw[1][2]),
    .valid_o_cast_nw                (valid_i_cast_nw[1][2]),
    .data_o_cast_nw                 (data_i_cast_nw[1][2]),
    .ready_i_cast_nw                (ready_o_cast_nw[1][2]),

    .valid_i_gather_nw              (valid_o_gather_nw[1][2]),
    .data_i_gather_nw               (data_o_gather_nw[1][2]),
    .ready_o_gather_nw              (ready_i_gather_nw[1][2]),
    .valid_o_gather_nw              (valid_i_gather_nw[1][2]),
    .data_o_gather_nw               (data_i_gather_nw[1][2]),
    .ready_i_gather_nw              (ready_o_gather_nw[1][2]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[1][2]),
    .data_i_merge_nw                (data_o_merge_nw[1][2]),
    .ready_o_merge_nw               (ready_i_merge_nw[1][2]),
    .valid_o_merge_nw               (valid_i_merge_nw[1][2]),
    .data_o_merge_nw                (data_i_merge_nw[1][2]),
    .ready_i_merge_nw               (ready_o_merge_nw[1][2]),

    .valid_i_cast_pe                (cast_valid_i_1_2),
    .data_i_cast_pe                 (cast_data_i_1_2),
    .ready_o_cast_pe                (cast_ready_o_1_2),
    .valid_o_cast_pe                (cast_valid_o_1_2),
    .data_o_cast_pe                 (cast_data_o_1_2),
    .ready_i_cast_pe                (cast_ready_i_1_2),

    .valid_i_merge_pe               (merge_valid_i_1_2),
    .data_i_merge_pe                (merge_data_i_1_2),
    .ready_o_merge_pe               (merge_ready_o_1_2),
    .valid_o_merge_pe               (merge_valid_o_1_2),
    .data_o_merge_pe                (merge_data_o_1_2),
    .ready_i_merge_pe               (merge_ready_i_1_2),

    .valid_i_gather_pe              (gather_valid_i_1_2),
    .data_i_gather_pe               (gather_data_i_1_2),
    .ready_o_gather_pe              (gather_ready_o_1_2),
    .valid_o_gather_pe              (gather_valid_o_1_2),
    .data_o_gather_pe               (gather_data_o_1_2),
    .ready_i_gather_pe              (gather_ready_i_1_2),

    .credit_upd                     (credit_upd[1][2])
);


network_interface #(
    .cast_out                       (cast_out_1_3),
    .gather_out                     (gather_out_1_3),
    .cast_sid                       (cast_sid_1_3),
    .gather_sid                     (gather_sid_1_3)
)ni_1_3(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[1][3]),
    .data_i_cast_nw                 (data_o_cast_nw[1][3]),
    .ready_o_cast_nw                (ready_i_cast_nw[1][3]),
    .valid_o_cast_nw                (valid_i_cast_nw[1][3]),
    .data_o_cast_nw                 (data_i_cast_nw[1][3]),
    .ready_i_cast_nw                (ready_o_cast_nw[1][3]),

    .valid_i_gather_nw              (valid_o_gather_nw[1][3]),
    .data_i_gather_nw               (data_o_gather_nw[1][3]),
    .ready_o_gather_nw              (ready_i_gather_nw[1][3]),
    .valid_o_gather_nw              (valid_i_gather_nw[1][3]),
    .data_o_gather_nw               (data_i_gather_nw[1][3]),
    .ready_i_gather_nw              (ready_o_gather_nw[1][3]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[1][3]),
    .data_i_merge_nw                (data_o_merge_nw[1][3]),
    .ready_o_merge_nw               (ready_i_merge_nw[1][3]),
    .valid_o_merge_nw               (valid_i_merge_nw[1][3]),
    .data_o_merge_nw                (data_i_merge_nw[1][3]),
    .ready_i_merge_nw               (ready_o_merge_nw[1][3]),

    .valid_i_cast_pe                (cast_valid_i_1_3),
    .data_i_cast_pe                 (cast_data_i_1_3),
    .ready_o_cast_pe                (cast_ready_o_1_3),
    .valid_o_cast_pe                (cast_valid_o_1_3),
    .data_o_cast_pe                 (cast_data_o_1_3),
    .ready_i_cast_pe                (cast_ready_i_1_3),

    .valid_i_merge_pe               (merge_valid_i_1_3),
    .data_i_merge_pe                (merge_data_i_1_3),
    .ready_o_merge_pe               (merge_ready_o_1_3),
    .valid_o_merge_pe               (merge_valid_o_1_3),
    .data_o_merge_pe                (merge_data_o_1_3),
    .ready_i_merge_pe               (merge_ready_i_1_3),

    .valid_i_gather_pe              (gather_valid_i_1_3),
    .data_i_gather_pe               (gather_data_i_1_3),
    .ready_o_gather_pe              (gather_ready_o_1_3),
    .valid_o_gather_pe              (gather_valid_o_1_3),
    .data_o_gather_pe               (gather_data_o_1_3),
    .ready_i_gather_pe              (gather_ready_i_1_3),

    .credit_upd                     (credit_upd[1][3])
);


network_interface #(
    .cast_out                       (cast_out_1_4),
    .gather_out                     (gather_out_1_4),
    .cast_sid                       (cast_sid_1_4),
    .gather_sid                     (gather_sid_1_4)
)ni_1_4(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[1][4]),
    .data_i_cast_nw                 (data_o_cast_nw[1][4]),
    .ready_o_cast_nw                (ready_i_cast_nw[1][4]),
    .valid_o_cast_nw                (valid_i_cast_nw[1][4]),
    .data_o_cast_nw                 (data_i_cast_nw[1][4]),
    .ready_i_cast_nw                (ready_o_cast_nw[1][4]),

    .valid_i_gather_nw              (valid_o_gather_nw[1][4]),
    .data_i_gather_nw               (data_o_gather_nw[1][4]),
    .ready_o_gather_nw              (ready_i_gather_nw[1][4]),
    .valid_o_gather_nw              (valid_i_gather_nw[1][4]),
    .data_o_gather_nw               (data_i_gather_nw[1][4]),
    .ready_i_gather_nw              (ready_o_gather_nw[1][4]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[1][4]),
    .data_i_merge_nw                (data_o_merge_nw[1][4]),
    .ready_o_merge_nw               (ready_i_merge_nw[1][4]),
    .valid_o_merge_nw               (valid_i_merge_nw[1][4]),
    .data_o_merge_nw                (data_i_merge_nw[1][4]),
    .ready_i_merge_nw               (ready_o_merge_nw[1][4]),

    .valid_i_cast_pe                (cast_valid_i_1_4),
    .data_i_cast_pe                 (cast_data_i_1_4),
    .ready_o_cast_pe                (cast_ready_o_1_4),
    .valid_o_cast_pe                (cast_valid_o_1_4),
    .data_o_cast_pe                 (cast_data_o_1_4),
    .ready_i_cast_pe                (cast_ready_i_1_4),

    .valid_i_merge_pe               (merge_valid_i_1_4),
    .data_i_merge_pe                (merge_data_i_1_4),
    .ready_o_merge_pe               (merge_ready_o_1_4),
    .valid_o_merge_pe               (merge_valid_o_1_4),
    .data_o_merge_pe                (merge_data_o_1_4),
    .ready_i_merge_pe               (merge_ready_i_1_4),

    .valid_i_gather_pe              (gather_valid_i_1_4),
    .data_i_gather_pe               (gather_data_i_1_4),
    .ready_o_gather_pe              (gather_ready_o_1_4),
    .valid_o_gather_pe              (gather_valid_o_1_4),
    .data_o_gather_pe               (gather_data_o_1_4),
    .ready_i_gather_pe              (gather_ready_i_1_4),

    .credit_upd                     (credit_upd[1][4])
);


network_interface #(
    .cast_out                       (cast_out_1_5),
    .gather_out                     (gather_out_1_5),
    .cast_sid                       (cast_sid_1_5),
    .gather_sid                     (gather_sid_1_5)
)ni_1_5(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[1][5]),
    .data_i_cast_nw                 (data_o_cast_nw[1][5]),
    .ready_o_cast_nw                (ready_i_cast_nw[1][5]),
    .valid_o_cast_nw                (valid_i_cast_nw[1][5]),
    .data_o_cast_nw                 (data_i_cast_nw[1][5]),
    .ready_i_cast_nw                (ready_o_cast_nw[1][5]),

    .valid_i_gather_nw              (valid_o_gather_nw[1][5]),
    .data_i_gather_nw               (data_o_gather_nw[1][5]),
    .ready_o_gather_nw              (ready_i_gather_nw[1][5]),
    .valid_o_gather_nw              (valid_i_gather_nw[1][5]),
    .data_o_gather_nw               (data_i_gather_nw[1][5]),
    .ready_i_gather_nw              (ready_o_gather_nw[1][5]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[1][5]),
    .data_i_merge_nw                (data_o_merge_nw[1][5]),
    .ready_o_merge_nw               (ready_i_merge_nw[1][5]),
    .valid_o_merge_nw               (valid_i_merge_nw[1][5]),
    .data_o_merge_nw                (data_i_merge_nw[1][5]),
    .ready_i_merge_nw               (ready_o_merge_nw[1][5]),

    .valid_i_cast_pe                (cast_valid_i_1_5),
    .data_i_cast_pe                 (cast_data_i_1_5),
    .ready_o_cast_pe                (cast_ready_o_1_5),
    .valid_o_cast_pe                (cast_valid_o_1_5),
    .data_o_cast_pe                 (cast_data_o_1_5),
    .ready_i_cast_pe                (cast_ready_i_1_5),

    .valid_i_merge_pe               (merge_valid_i_1_5),
    .data_i_merge_pe                (merge_data_i_1_5),
    .ready_o_merge_pe               (merge_ready_o_1_5),
    .valid_o_merge_pe               (merge_valid_o_1_5),
    .data_o_merge_pe                (merge_data_o_1_5),
    .ready_i_merge_pe               (merge_ready_i_1_5),

    .valid_i_gather_pe              (gather_valid_i_1_5),
    .data_i_gather_pe               (gather_data_i_1_5),
    .ready_o_gather_pe              (gather_ready_o_1_5),
    .valid_o_gather_pe              (gather_valid_o_1_5),
    .data_o_gather_pe               (gather_data_o_1_5),
    .ready_i_gather_pe              (gather_ready_i_1_5),

    .credit_upd                     (credit_upd[1][5])
);


network_interface #(
    .cast_out                       (cast_out_1_6),
    .gather_out                     (gather_out_1_6),
    .cast_sid                       (cast_sid_1_6),
    .gather_sid                     (gather_sid_1_6)
)ni_1_6(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[1][6]),
    .data_i_cast_nw                 (data_o_cast_nw[1][6]),
    .ready_o_cast_nw                (ready_i_cast_nw[1][6]),
    .valid_o_cast_nw                (valid_i_cast_nw[1][6]),
    .data_o_cast_nw                 (data_i_cast_nw[1][6]),
    .ready_i_cast_nw                (ready_o_cast_nw[1][6]),

    .valid_i_gather_nw              (valid_o_gather_nw[1][6]),
    .data_i_gather_nw               (data_o_gather_nw[1][6]),
    .ready_o_gather_nw              (ready_i_gather_nw[1][6]),
    .valid_o_gather_nw              (valid_i_gather_nw[1][6]),
    .data_o_gather_nw               (data_i_gather_nw[1][6]),
    .ready_i_gather_nw              (ready_o_gather_nw[1][6]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[1][6]),
    .data_i_merge_nw                (data_o_merge_nw[1][6]),
    .ready_o_merge_nw               (ready_i_merge_nw[1][6]),
    .valid_o_merge_nw               (valid_i_merge_nw[1][6]),
    .data_o_merge_nw                (data_i_merge_nw[1][6]),
    .ready_i_merge_nw               (ready_o_merge_nw[1][6]),

    .valid_i_cast_pe                (cast_valid_i_1_6),
    .data_i_cast_pe                 (cast_data_i_1_6),
    .ready_o_cast_pe                (cast_ready_o_1_6),
    .valid_o_cast_pe                (cast_valid_o_1_6),
    .data_o_cast_pe                 (cast_data_o_1_6),
    .ready_i_cast_pe                (cast_ready_i_1_6),

    .valid_i_merge_pe               (merge_valid_i_1_6),
    .data_i_merge_pe                (merge_data_i_1_6),
    .ready_o_merge_pe               (merge_ready_o_1_6),
    .valid_o_merge_pe               (merge_valid_o_1_6),
    .data_o_merge_pe                (merge_data_o_1_6),
    .ready_i_merge_pe               (merge_ready_i_1_6),

    .valid_i_gather_pe              (gather_valid_i_1_6),
    .data_i_gather_pe               (gather_data_i_1_6),
    .ready_o_gather_pe              (gather_ready_o_1_6),
    .valid_o_gather_pe              (gather_valid_o_1_6),
    .data_o_gather_pe               (gather_data_o_1_6),
    .ready_i_gather_pe              (gather_ready_i_1_6),

    .credit_upd                     (credit_upd[1][6])
);


network_interface #(
    .cast_out                       (cast_out_1_7),
    .gather_out                     (gather_out_1_7),
    .cast_sid                       (cast_sid_1_7),
    .gather_sid                     (gather_sid_1_7)
)ni_1_7(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[1][7]),
    .data_i_cast_nw                 (data_o_cast_nw[1][7]),
    .ready_o_cast_nw                (ready_i_cast_nw[1][7]),
    .valid_o_cast_nw                (valid_i_cast_nw[1][7]),
    .data_o_cast_nw                 (data_i_cast_nw[1][7]),
    .ready_i_cast_nw                (ready_o_cast_nw[1][7]),

    .valid_i_gather_nw              (valid_o_gather_nw[1][7]),
    .data_i_gather_nw               (data_o_gather_nw[1][7]),
    .ready_o_gather_nw              (ready_i_gather_nw[1][7]),
    .valid_o_gather_nw              (valid_i_gather_nw[1][7]),
    .data_o_gather_nw               (data_i_gather_nw[1][7]),
    .ready_i_gather_nw              (ready_o_gather_nw[1][7]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[1][7]),
    .data_i_merge_nw                (data_o_merge_nw[1][7]),
    .ready_o_merge_nw               (ready_i_merge_nw[1][7]),
    .valid_o_merge_nw               (valid_i_merge_nw[1][7]),
    .data_o_merge_nw                (data_i_merge_nw[1][7]),
    .ready_i_merge_nw               (ready_o_merge_nw[1][7]),

    .valid_i_cast_pe                (cast_valid_i_1_7),
    .data_i_cast_pe                 (cast_data_i_1_7),
    .ready_o_cast_pe                (cast_ready_o_1_7),
    .valid_o_cast_pe                (cast_valid_o_1_7),
    .data_o_cast_pe                 (cast_data_o_1_7),
    .ready_i_cast_pe                (cast_ready_i_1_7),

    .valid_i_merge_pe               (merge_valid_i_1_7),
    .data_i_merge_pe                (merge_data_i_1_7),
    .ready_o_merge_pe               (merge_ready_o_1_7),
    .valid_o_merge_pe               (merge_valid_o_1_7),
    .data_o_merge_pe                (merge_data_o_1_7),
    .ready_i_merge_pe               (merge_ready_i_1_7),

    .valid_i_gather_pe              (gather_valid_i_1_7),
    .data_i_gather_pe               (gather_data_i_1_7),
    .ready_o_gather_pe              (gather_ready_o_1_7),
    .valid_o_gather_pe              (gather_valid_o_1_7),
    .data_o_gather_pe               (gather_data_o_1_7),
    .ready_i_gather_pe              (gather_ready_i_1_7),

    .credit_upd                     (credit_upd[1][7])
);


network_interface #(
    .cast_out                       (cast_out_1_8),
    .gather_out                     (gather_out_1_8),
    .cast_sid                       (cast_sid_1_8),
    .gather_sid                     (gather_sid_1_8)
)ni_1_8(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[1][8]),
    .data_i_cast_nw                 (data_o_cast_nw[1][8]),
    .ready_o_cast_nw                (ready_i_cast_nw[1][8]),
    .valid_o_cast_nw                (valid_i_cast_nw[1][8]),
    .data_o_cast_nw                 (data_i_cast_nw[1][8]),
    .ready_i_cast_nw                (ready_o_cast_nw[1][8]),

    .valid_i_gather_nw              (valid_o_gather_nw[1][8]),
    .data_i_gather_nw               (data_o_gather_nw[1][8]),
    .ready_o_gather_nw              (ready_i_gather_nw[1][8]),
    .valid_o_gather_nw              (valid_i_gather_nw[1][8]),
    .data_o_gather_nw               (data_i_gather_nw[1][8]),
    .ready_i_gather_nw              (ready_o_gather_nw[1][8]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[1][8]),
    .data_i_merge_nw                (data_o_merge_nw[1][8]),
    .ready_o_merge_nw               (ready_i_merge_nw[1][8]),
    .valid_o_merge_nw               (valid_i_merge_nw[1][8]),
    .data_o_merge_nw                (data_i_merge_nw[1][8]),
    .ready_i_merge_nw               (ready_o_merge_nw[1][8]),

    .valid_i_cast_pe                (cast_valid_i_1_8),
    .data_i_cast_pe                 (cast_data_i_1_8),
    .ready_o_cast_pe                (cast_ready_o_1_8),
    .valid_o_cast_pe                (cast_valid_o_1_8),
    .data_o_cast_pe                 (cast_data_o_1_8),
    .ready_i_cast_pe                (cast_ready_i_1_8),

    .valid_i_merge_pe               (merge_valid_i_1_8),
    .data_i_merge_pe                (merge_data_i_1_8),
    .ready_o_merge_pe               (merge_ready_o_1_8),
    .valid_o_merge_pe               (merge_valid_o_1_8),
    .data_o_merge_pe                (merge_data_o_1_8),
    .ready_i_merge_pe               (merge_ready_i_1_8),

    .valid_i_gather_pe              (gather_valid_i_1_8),
    .data_i_gather_pe               (gather_data_i_1_8),
    .ready_o_gather_pe              (gather_ready_o_1_8),
    .valid_o_gather_pe              (gather_valid_o_1_8),
    .data_o_gather_pe               (gather_data_o_1_8),
    .ready_i_gather_pe              (gather_ready_i_1_8),

    .credit_upd                     (credit_upd[1][8])
);


network_interface #(
    .cast_out                       (cast_out_1_9),
    .gather_out                     (gather_out_1_9),
    .cast_sid                       (cast_sid_1_9),
    .gather_sid                     (gather_sid_1_9)
)ni_1_9(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[1][9]),
    .data_i_cast_nw                 (data_o_cast_nw[1][9]),
    .ready_o_cast_nw                (ready_i_cast_nw[1][9]),
    .valid_o_cast_nw                (valid_i_cast_nw[1][9]),
    .data_o_cast_nw                 (data_i_cast_nw[1][9]),
    .ready_i_cast_nw                (ready_o_cast_nw[1][9]),

    .valid_i_gather_nw              (valid_o_gather_nw[1][9]),
    .data_i_gather_nw               (data_o_gather_nw[1][9]),
    .ready_o_gather_nw              (ready_i_gather_nw[1][9]),
    .valid_o_gather_nw              (valid_i_gather_nw[1][9]),
    .data_o_gather_nw               (data_i_gather_nw[1][9]),
    .ready_i_gather_nw              (ready_o_gather_nw[1][9]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[1][9]),
    .data_i_merge_nw                (data_o_merge_nw[1][9]),
    .ready_o_merge_nw               (ready_i_merge_nw[1][9]),
    .valid_o_merge_nw               (valid_i_merge_nw[1][9]),
    .data_o_merge_nw                (data_i_merge_nw[1][9]),
    .ready_i_merge_nw               (ready_o_merge_nw[1][9]),

    .valid_i_cast_pe                (cast_valid_i_1_9),
    .data_i_cast_pe                 (cast_data_i_1_9),
    .ready_o_cast_pe                (cast_ready_o_1_9),
    .valid_o_cast_pe                (cast_valid_o_1_9),
    .data_o_cast_pe                 (cast_data_o_1_9),
    .ready_i_cast_pe                (cast_ready_i_1_9),

    .valid_i_merge_pe               (merge_valid_i_1_9),
    .data_i_merge_pe                (merge_data_i_1_9),
    .ready_o_merge_pe               (merge_ready_o_1_9),
    .valid_o_merge_pe               (merge_valid_o_1_9),
    .data_o_merge_pe                (merge_data_o_1_9),
    .ready_i_merge_pe               (merge_ready_i_1_9),

    .valid_i_gather_pe              (gather_valid_i_1_9),
    .data_i_gather_pe               (gather_data_i_1_9),
    .ready_o_gather_pe              (gather_ready_o_1_9),
    .valid_o_gather_pe              (gather_valid_o_1_9),
    .data_o_gather_pe               (gather_data_o_1_9),
    .ready_i_gather_pe              (gather_ready_i_1_9),

    .credit_upd                     (credit_upd[1][9])
);


network_interface #(
    .cast_out                       (cast_out_1_10),
    .gather_out                     (gather_out_1_10),
    .cast_sid                       (cast_sid_1_10),
    .gather_sid                     (gather_sid_1_10)
)ni_1_10(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[1][10]),
    .data_i_cast_nw                 (data_o_cast_nw[1][10]),
    .ready_o_cast_nw                (ready_i_cast_nw[1][10]),
    .valid_o_cast_nw                (valid_i_cast_nw[1][10]),
    .data_o_cast_nw                 (data_i_cast_nw[1][10]),
    .ready_i_cast_nw                (ready_o_cast_nw[1][10]),

    .valid_i_gather_nw              (valid_o_gather_nw[1][10]),
    .data_i_gather_nw               (data_o_gather_nw[1][10]),
    .ready_o_gather_nw              (ready_i_gather_nw[1][10]),
    .valid_o_gather_nw              (valid_i_gather_nw[1][10]),
    .data_o_gather_nw               (data_i_gather_nw[1][10]),
    .ready_i_gather_nw              (ready_o_gather_nw[1][10]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[1][10]),
    .data_i_merge_nw                (data_o_merge_nw[1][10]),
    .ready_o_merge_nw               (ready_i_merge_nw[1][10]),
    .valid_o_merge_nw               (valid_i_merge_nw[1][10]),
    .data_o_merge_nw                (data_i_merge_nw[1][10]),
    .ready_i_merge_nw               (ready_o_merge_nw[1][10]),

    .valid_i_cast_pe                (cast_valid_i_1_10),
    .data_i_cast_pe                 (cast_data_i_1_10),
    .ready_o_cast_pe                (cast_ready_o_1_10),
    .valid_o_cast_pe                (cast_valid_o_1_10),
    .data_o_cast_pe                 (cast_data_o_1_10),
    .ready_i_cast_pe                (cast_ready_i_1_10),

    .valid_i_merge_pe               (merge_valid_i_1_10),
    .data_i_merge_pe                (merge_data_i_1_10),
    .ready_o_merge_pe               (merge_ready_o_1_10),
    .valid_o_merge_pe               (merge_valid_o_1_10),
    .data_o_merge_pe                (merge_data_o_1_10),
    .ready_i_merge_pe               (merge_ready_i_1_10),

    .valid_i_gather_pe              (gather_valid_i_1_10),
    .data_i_gather_pe               (gather_data_i_1_10),
    .ready_o_gather_pe              (gather_ready_o_1_10),
    .valid_o_gather_pe              (gather_valid_o_1_10),
    .data_o_gather_pe               (gather_data_o_1_10),
    .ready_i_gather_pe              (gather_ready_i_1_10),

    .credit_upd                     (credit_upd[1][10])
);


network_interface #(
    .cast_out                       (cast_out_1_11),
    .gather_out                     (gather_out_1_11),
    .cast_sid                       (cast_sid_1_11),
    .gather_sid                     (gather_sid_1_11)
)ni_1_11(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[1][11]),
    .data_i_cast_nw                 (data_o_cast_nw[1][11]),
    .ready_o_cast_nw                (ready_i_cast_nw[1][11]),
    .valid_o_cast_nw                (valid_i_cast_nw[1][11]),
    .data_o_cast_nw                 (data_i_cast_nw[1][11]),
    .ready_i_cast_nw                (ready_o_cast_nw[1][11]),

    .valid_i_gather_nw              (valid_o_gather_nw[1][11]),
    .data_i_gather_nw               (data_o_gather_nw[1][11]),
    .ready_o_gather_nw              (ready_i_gather_nw[1][11]),
    .valid_o_gather_nw              (valid_i_gather_nw[1][11]),
    .data_o_gather_nw               (data_i_gather_nw[1][11]),
    .ready_i_gather_nw              (ready_o_gather_nw[1][11]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[1][11]),
    .data_i_merge_nw                (data_o_merge_nw[1][11]),
    .ready_o_merge_nw               (ready_i_merge_nw[1][11]),
    .valid_o_merge_nw               (valid_i_merge_nw[1][11]),
    .data_o_merge_nw                (data_i_merge_nw[1][11]),
    .ready_i_merge_nw               (ready_o_merge_nw[1][11]),

    .valid_i_cast_pe                (cast_valid_i_1_11),
    .data_i_cast_pe                 (cast_data_i_1_11),
    .ready_o_cast_pe                (cast_ready_o_1_11),
    .valid_o_cast_pe                (cast_valid_o_1_11),
    .data_o_cast_pe                 (cast_data_o_1_11),
    .ready_i_cast_pe                (cast_ready_i_1_11),

    .valid_i_merge_pe               (merge_valid_i_1_11),
    .data_i_merge_pe                (merge_data_i_1_11),
    .ready_o_merge_pe               (merge_ready_o_1_11),
    .valid_o_merge_pe               (merge_valid_o_1_11),
    .data_o_merge_pe                (merge_data_o_1_11),
    .ready_i_merge_pe               (merge_ready_i_1_11),

    .valid_i_gather_pe              (gather_valid_i_1_11),
    .data_i_gather_pe               (gather_data_i_1_11),
    .ready_o_gather_pe              (gather_ready_o_1_11),
    .valid_o_gather_pe              (gather_valid_o_1_11),
    .data_o_gather_pe               (gather_data_o_1_11),
    .ready_i_gather_pe              (gather_ready_i_1_11),

    .credit_upd                     (credit_upd[1][11])
);


network_interface #(
    .cast_out                       (cast_out_1_12),
    .gather_out                     (gather_out_1_12),
    .cast_sid                       (cast_sid_1_12),
    .gather_sid                     (gather_sid_1_12)
)ni_1_12(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[1][12]),
    .data_i_cast_nw                 (data_o_cast_nw[1][12]),
    .ready_o_cast_nw                (ready_i_cast_nw[1][12]),
    .valid_o_cast_nw                (valid_i_cast_nw[1][12]),
    .data_o_cast_nw                 (data_i_cast_nw[1][12]),
    .ready_i_cast_nw                (ready_o_cast_nw[1][12]),

    .valid_i_gather_nw              (valid_o_gather_nw[1][12]),
    .data_i_gather_nw               (data_o_gather_nw[1][12]),
    .ready_o_gather_nw              (ready_i_gather_nw[1][12]),
    .valid_o_gather_nw              (valid_i_gather_nw[1][12]),
    .data_o_gather_nw               (data_i_gather_nw[1][12]),
    .ready_i_gather_nw              (ready_o_gather_nw[1][12]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[1][12]),
    .data_i_merge_nw                (data_o_merge_nw[1][12]),
    .ready_o_merge_nw               (ready_i_merge_nw[1][12]),
    .valid_o_merge_nw               (valid_i_merge_nw[1][12]),
    .data_o_merge_nw                (data_i_merge_nw[1][12]),
    .ready_i_merge_nw               (ready_o_merge_nw[1][12]),

    .valid_i_cast_pe                (cast_valid_i_1_12),
    .data_i_cast_pe                 (cast_data_i_1_12),
    .ready_o_cast_pe                (cast_ready_o_1_12),
    .valid_o_cast_pe                (cast_valid_o_1_12),
    .data_o_cast_pe                 (cast_data_o_1_12),
    .ready_i_cast_pe                (cast_ready_i_1_12),

    .valid_i_merge_pe               (merge_valid_i_1_12),
    .data_i_merge_pe                (merge_data_i_1_12),
    .ready_o_merge_pe               (merge_ready_o_1_12),
    .valid_o_merge_pe               (merge_valid_o_1_12),
    .data_o_merge_pe                (merge_data_o_1_12),
    .ready_i_merge_pe               (merge_ready_i_1_12),

    .valid_i_gather_pe              (gather_valid_i_1_12),
    .data_i_gather_pe               (gather_data_i_1_12),
    .ready_o_gather_pe              (gather_ready_o_1_12),
    .valid_o_gather_pe              (gather_valid_o_1_12),
    .data_o_gather_pe               (gather_data_o_1_12),
    .ready_i_gather_pe              (gather_ready_i_1_12),

    .credit_upd                     (credit_upd[1][12])
);


network_interface #(
    .cast_out                       (cast_out_1_13),
    .gather_out                     (gather_out_1_13),
    .cast_sid                       (cast_sid_1_13),
    .gather_sid                     (gather_sid_1_13)
)ni_1_13(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[1][13]),
    .data_i_cast_nw                 (data_o_cast_nw[1][13]),
    .ready_o_cast_nw                (ready_i_cast_nw[1][13]),
    .valid_o_cast_nw                (valid_i_cast_nw[1][13]),
    .data_o_cast_nw                 (data_i_cast_nw[1][13]),
    .ready_i_cast_nw                (ready_o_cast_nw[1][13]),

    .valid_i_gather_nw              (valid_o_gather_nw[1][13]),
    .data_i_gather_nw               (data_o_gather_nw[1][13]),
    .ready_o_gather_nw              (ready_i_gather_nw[1][13]),
    .valid_o_gather_nw              (valid_i_gather_nw[1][13]),
    .data_o_gather_nw               (data_i_gather_nw[1][13]),
    .ready_i_gather_nw              (ready_o_gather_nw[1][13]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[1][13]),
    .data_i_merge_nw                (data_o_merge_nw[1][13]),
    .ready_o_merge_nw               (ready_i_merge_nw[1][13]),
    .valid_o_merge_nw               (valid_i_merge_nw[1][13]),
    .data_o_merge_nw                (data_i_merge_nw[1][13]),
    .ready_i_merge_nw               (ready_o_merge_nw[1][13]),

    .valid_i_cast_pe                (cast_valid_i_1_13),
    .data_i_cast_pe                 (cast_data_i_1_13),
    .ready_o_cast_pe                (cast_ready_o_1_13),
    .valid_o_cast_pe                (cast_valid_o_1_13),
    .data_o_cast_pe                 (cast_data_o_1_13),
    .ready_i_cast_pe                (cast_ready_i_1_13),

    .valid_i_merge_pe               (merge_valid_i_1_13),
    .data_i_merge_pe                (merge_data_i_1_13),
    .ready_o_merge_pe               (merge_ready_o_1_13),
    .valid_o_merge_pe               (merge_valid_o_1_13),
    .data_o_merge_pe                (merge_data_o_1_13),
    .ready_i_merge_pe               (merge_ready_i_1_13),

    .valid_i_gather_pe              (gather_valid_i_1_13),
    .data_i_gather_pe               (gather_data_i_1_13),
    .ready_o_gather_pe              (gather_ready_o_1_13),
    .valid_o_gather_pe              (gather_valid_o_1_13),
    .data_o_gather_pe               (gather_data_o_1_13),
    .ready_i_gather_pe              (gather_ready_i_1_13),

    .credit_upd                     (credit_upd[1][13])
);


network_interface #(
    .cast_out                       (cast_out_1_14),
    .gather_out                     (gather_out_1_14),
    .cast_sid                       (cast_sid_1_14),
    .gather_sid                     (gather_sid_1_14)
)ni_1_14(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[1][14]),
    .data_i_cast_nw                 (data_o_cast_nw[1][14]),
    .ready_o_cast_nw                (ready_i_cast_nw[1][14]),
    .valid_o_cast_nw                (valid_i_cast_nw[1][14]),
    .data_o_cast_nw                 (data_i_cast_nw[1][14]),
    .ready_i_cast_nw                (ready_o_cast_nw[1][14]),

    .valid_i_gather_nw              (valid_o_gather_nw[1][14]),
    .data_i_gather_nw               (data_o_gather_nw[1][14]),
    .ready_o_gather_nw              (ready_i_gather_nw[1][14]),
    .valid_o_gather_nw              (valid_i_gather_nw[1][14]),
    .data_o_gather_nw               (data_i_gather_nw[1][14]),
    .ready_i_gather_nw              (ready_o_gather_nw[1][14]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[1][14]),
    .data_i_merge_nw                (data_o_merge_nw[1][14]),
    .ready_o_merge_nw               (ready_i_merge_nw[1][14]),
    .valid_o_merge_nw               (valid_i_merge_nw[1][14]),
    .data_o_merge_nw                (data_i_merge_nw[1][14]),
    .ready_i_merge_nw               (ready_o_merge_nw[1][14]),

    .valid_i_cast_pe                (cast_valid_i_1_14),
    .data_i_cast_pe                 (cast_data_i_1_14),
    .ready_o_cast_pe                (cast_ready_o_1_14),
    .valid_o_cast_pe                (cast_valid_o_1_14),
    .data_o_cast_pe                 (cast_data_o_1_14),
    .ready_i_cast_pe                (cast_ready_i_1_14),

    .valid_i_merge_pe               (merge_valid_i_1_14),
    .data_i_merge_pe                (merge_data_i_1_14),
    .ready_o_merge_pe               (merge_ready_o_1_14),
    .valid_o_merge_pe               (merge_valid_o_1_14),
    .data_o_merge_pe                (merge_data_o_1_14),
    .ready_i_merge_pe               (merge_ready_i_1_14),

    .valid_i_gather_pe              (gather_valid_i_1_14),
    .data_i_gather_pe               (gather_data_i_1_14),
    .ready_o_gather_pe              (gather_ready_o_1_14),
    .valid_o_gather_pe              (gather_valid_o_1_14),
    .data_o_gather_pe               (gather_data_o_1_14),
    .ready_i_gather_pe              (gather_ready_i_1_14),

    .credit_upd                     (credit_upd[1][14])
);


network_interface #(
    .cast_out                       (cast_out_1_15),
    .gather_out                     (gather_out_1_15),
    .cast_sid                       (cast_sid_1_15),
    .gather_sid                     (gather_sid_1_15)
)ni_1_15(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[1][15]),
    .data_i_cast_nw                 (data_o_cast_nw[1][15]),
    .ready_o_cast_nw                (ready_i_cast_nw[1][15]),
    .valid_o_cast_nw                (valid_i_cast_nw[1][15]),
    .data_o_cast_nw                 (data_i_cast_nw[1][15]),
    .ready_i_cast_nw                (ready_o_cast_nw[1][15]),

    .valid_i_gather_nw              (valid_o_gather_nw[1][15]),
    .data_i_gather_nw               (data_o_gather_nw[1][15]),
    .ready_o_gather_nw              (ready_i_gather_nw[1][15]),
    .valid_o_gather_nw              (valid_i_gather_nw[1][15]),
    .data_o_gather_nw               (data_i_gather_nw[1][15]),
    .ready_i_gather_nw              (ready_o_gather_nw[1][15]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[1][15]),
    .data_i_merge_nw                (data_o_merge_nw[1][15]),
    .ready_o_merge_nw               (ready_i_merge_nw[1][15]),
    .valid_o_merge_nw               (valid_i_merge_nw[1][15]),
    .data_o_merge_nw                (data_i_merge_nw[1][15]),
    .ready_i_merge_nw               (ready_o_merge_nw[1][15]),

    .valid_i_cast_pe                (cast_valid_i_1_15),
    .data_i_cast_pe                 (cast_data_i_1_15),
    .ready_o_cast_pe                (cast_ready_o_1_15),
    .valid_o_cast_pe                (cast_valid_o_1_15),
    .data_o_cast_pe                 (cast_data_o_1_15),
    .ready_i_cast_pe                (cast_ready_i_1_15),

    .valid_i_merge_pe               (merge_valid_i_1_15),
    .data_i_merge_pe                (merge_data_i_1_15),
    .ready_o_merge_pe               (merge_ready_o_1_15),
    .valid_o_merge_pe               (merge_valid_o_1_15),
    .data_o_merge_pe                (merge_data_o_1_15),
    .ready_i_merge_pe               (merge_ready_i_1_15),

    .valid_i_gather_pe              (gather_valid_i_1_15),
    .data_i_gather_pe               (gather_data_i_1_15),
    .ready_o_gather_pe              (gather_ready_o_1_15),
    .valid_o_gather_pe              (gather_valid_o_1_15),
    .data_o_gather_pe               (gather_data_o_1_15),
    .ready_i_gather_pe              (gather_ready_i_1_15),

    .credit_upd                     (credit_upd[1][15])
);


network_interface #(
    .cast_out                       (cast_out_1_16),
    .gather_out                     (gather_out_1_16),
    .cast_sid                       (cast_sid_1_16),
    .gather_sid                     (gather_sid_1_16)
)ni_1_16(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[1][16]),
    .data_i_cast_nw                 (data_o_cast_nw[1][16]),
    .ready_o_cast_nw                (ready_i_cast_nw[1][16]),
    .valid_o_cast_nw                (valid_i_cast_nw[1][16]),
    .data_o_cast_nw                 (data_i_cast_nw[1][16]),
    .ready_i_cast_nw                (ready_o_cast_nw[1][16]),

    .valid_i_gather_nw              (valid_o_gather_nw[1][16]),
    .data_i_gather_nw               (data_o_gather_nw[1][16]),
    .ready_o_gather_nw              (ready_i_gather_nw[1][16]),
    .valid_o_gather_nw              (valid_i_gather_nw[1][16]),
    .data_o_gather_nw               (data_i_gather_nw[1][16]),
    .ready_i_gather_nw              (ready_o_gather_nw[1][16]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[1][16]),
    .data_i_merge_nw                (data_o_merge_nw[1][16]),
    .ready_o_merge_nw               (ready_i_merge_nw[1][16]),
    .valid_o_merge_nw               (valid_i_merge_nw[1][16]),
    .data_o_merge_nw                (data_i_merge_nw[1][16]),
    .ready_i_merge_nw               (ready_o_merge_nw[1][16]),

    .valid_i_cast_pe                (cast_valid_i_1_16),
    .data_i_cast_pe                 (cast_data_i_1_16),
    .ready_o_cast_pe                (cast_ready_o_1_16),
    .valid_o_cast_pe                (cast_valid_o_1_16),
    .data_o_cast_pe                 (cast_data_o_1_16),
    .ready_i_cast_pe                (cast_ready_i_1_16),

    .valid_i_merge_pe               (merge_valid_i_1_16),
    .data_i_merge_pe                (merge_data_i_1_16),
    .ready_o_merge_pe               (merge_ready_o_1_16),
    .valid_o_merge_pe               (merge_valid_o_1_16),
    .data_o_merge_pe                (merge_data_o_1_16),
    .ready_i_merge_pe               (merge_ready_i_1_16),

    .valid_i_gather_pe              (gather_valid_i_1_16),
    .data_i_gather_pe               (gather_data_i_1_16),
    .ready_o_gather_pe              (gather_ready_o_1_16),
    .valid_o_gather_pe              (gather_valid_o_1_16),
    .data_o_gather_pe               (gather_data_o_1_16),
    .ready_i_gather_pe              (gather_ready_i_1_16),

    .credit_upd                     (credit_upd[1][16])
);


network_interface #(
    .cast_out                       (cast_out_1_17),
    .gather_out                     (gather_out_1_17),
    .cast_sid                       (cast_sid_1_17),
    .gather_sid                     (gather_sid_1_17)
)ni_1_17(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[1][17]),
    .data_i_cast_nw                 (data_o_cast_nw[1][17]),
    .ready_o_cast_nw                (ready_i_cast_nw[1][17]),
    .valid_o_cast_nw                (valid_i_cast_nw[1][17]),
    .data_o_cast_nw                 (data_i_cast_nw[1][17]),
    .ready_i_cast_nw                (ready_o_cast_nw[1][17]),

    .valid_i_gather_nw              (valid_o_gather_nw[1][17]),
    .data_i_gather_nw               (data_o_gather_nw[1][17]),
    .ready_o_gather_nw              (ready_i_gather_nw[1][17]),
    .valid_o_gather_nw              (valid_i_gather_nw[1][17]),
    .data_o_gather_nw               (data_i_gather_nw[1][17]),
    .ready_i_gather_nw              (ready_o_gather_nw[1][17]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[1][17]),
    .data_i_merge_nw                (data_o_merge_nw[1][17]),
    .ready_o_merge_nw               (ready_i_merge_nw[1][17]),
    .valid_o_merge_nw               (valid_i_merge_nw[1][17]),
    .data_o_merge_nw                (data_i_merge_nw[1][17]),
    .ready_i_merge_nw               (ready_o_merge_nw[1][17]),

    .valid_i_cast_pe                (cast_valid_i_1_17),
    .data_i_cast_pe                 (cast_data_i_1_17),
    .ready_o_cast_pe                (cast_ready_o_1_17),
    .valid_o_cast_pe                (cast_valid_o_1_17),
    .data_o_cast_pe                 (cast_data_o_1_17),
    .ready_i_cast_pe                (cast_ready_i_1_17),

    .valid_i_merge_pe               (merge_valid_i_1_17),
    .data_i_merge_pe                (merge_data_i_1_17),
    .ready_o_merge_pe               (merge_ready_o_1_17),
    .valid_o_merge_pe               (merge_valid_o_1_17),
    .data_o_merge_pe                (merge_data_o_1_17),
    .ready_i_merge_pe               (merge_ready_i_1_17),

    .valid_i_gather_pe              (gather_valid_i_1_17),
    .data_i_gather_pe               (gather_data_i_1_17),
    .ready_o_gather_pe              (gather_ready_o_1_17),
    .valid_o_gather_pe              (gather_valid_o_1_17),
    .data_o_gather_pe               (gather_data_o_1_17),
    .ready_i_gather_pe              (gather_ready_i_1_17),

    .credit_upd                     (credit_upd[1][17])
);


network_interface #(
    .cast_out                       (cast_out_1_18),
    .gather_out                     (gather_out_1_18),
    .cast_sid                       (cast_sid_1_18),
    .gather_sid                     (gather_sid_1_18)
)ni_1_18(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[1][18]),
    .data_i_cast_nw                 (data_o_cast_nw[1][18]),
    .ready_o_cast_nw                (ready_i_cast_nw[1][18]),
    .valid_o_cast_nw                (valid_i_cast_nw[1][18]),
    .data_o_cast_nw                 (data_i_cast_nw[1][18]),
    .ready_i_cast_nw                (ready_o_cast_nw[1][18]),

    .valid_i_gather_nw              (valid_o_gather_nw[1][18]),
    .data_i_gather_nw               (data_o_gather_nw[1][18]),
    .ready_o_gather_nw              (ready_i_gather_nw[1][18]),
    .valid_o_gather_nw              (valid_i_gather_nw[1][18]),
    .data_o_gather_nw               (data_i_gather_nw[1][18]),
    .ready_i_gather_nw              (ready_o_gather_nw[1][18]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[1][18]),
    .data_i_merge_nw                (data_o_merge_nw[1][18]),
    .ready_o_merge_nw               (ready_i_merge_nw[1][18]),
    .valid_o_merge_nw               (valid_i_merge_nw[1][18]),
    .data_o_merge_nw                (data_i_merge_nw[1][18]),
    .ready_i_merge_nw               (ready_o_merge_nw[1][18]),

    .valid_i_cast_pe                (cast_valid_i_1_18),
    .data_i_cast_pe                 (cast_data_i_1_18),
    .ready_o_cast_pe                (cast_ready_o_1_18),
    .valid_o_cast_pe                (cast_valid_o_1_18),
    .data_o_cast_pe                 (cast_data_o_1_18),
    .ready_i_cast_pe                (cast_ready_i_1_18),

    .valid_i_merge_pe               (merge_valid_i_1_18),
    .data_i_merge_pe                (merge_data_i_1_18),
    .ready_o_merge_pe               (merge_ready_o_1_18),
    .valid_o_merge_pe               (merge_valid_o_1_18),
    .data_o_merge_pe                (merge_data_o_1_18),
    .ready_i_merge_pe               (merge_ready_i_1_18),

    .valid_i_gather_pe              (gather_valid_i_1_18),
    .data_i_gather_pe               (gather_data_i_1_18),
    .ready_o_gather_pe              (gather_ready_o_1_18),
    .valid_o_gather_pe              (gather_valid_o_1_18),
    .data_o_gather_pe               (gather_data_o_1_18),
    .ready_i_gather_pe              (gather_ready_i_1_18),

    .credit_upd                     (credit_upd[1][18])
);


network_interface #(
    .cast_out                       (cast_out_1_19),
    .gather_out                     (gather_out_1_19),
    .cast_sid                       (cast_sid_1_19),
    .gather_sid                     (gather_sid_1_19)
)ni_1_19(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[1][19]),
    .data_i_cast_nw                 (data_o_cast_nw[1][19]),
    .ready_o_cast_nw                (ready_i_cast_nw[1][19]),
    .valid_o_cast_nw                (valid_i_cast_nw[1][19]),
    .data_o_cast_nw                 (data_i_cast_nw[1][19]),
    .ready_i_cast_nw                (ready_o_cast_nw[1][19]),

    .valid_i_gather_nw              (valid_o_gather_nw[1][19]),
    .data_i_gather_nw               (data_o_gather_nw[1][19]),
    .ready_o_gather_nw              (ready_i_gather_nw[1][19]),
    .valid_o_gather_nw              (valid_i_gather_nw[1][19]),
    .data_o_gather_nw               (data_i_gather_nw[1][19]),
    .ready_i_gather_nw              (ready_o_gather_nw[1][19]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[1][19]),
    .data_i_merge_nw                (data_o_merge_nw[1][19]),
    .ready_o_merge_nw               (ready_i_merge_nw[1][19]),
    .valid_o_merge_nw               (valid_i_merge_nw[1][19]),
    .data_o_merge_nw                (data_i_merge_nw[1][19]),
    .ready_i_merge_nw               (ready_o_merge_nw[1][19]),

    .valid_i_cast_pe                (cast_valid_i_1_19),
    .data_i_cast_pe                 (cast_data_i_1_19),
    .ready_o_cast_pe                (cast_ready_o_1_19),
    .valid_o_cast_pe                (cast_valid_o_1_19),
    .data_o_cast_pe                 (cast_data_o_1_19),
    .ready_i_cast_pe                (cast_ready_i_1_19),

    .valid_i_merge_pe               (merge_valid_i_1_19),
    .data_i_merge_pe                (merge_data_i_1_19),
    .ready_o_merge_pe               (merge_ready_o_1_19),
    .valid_o_merge_pe               (merge_valid_o_1_19),
    .data_o_merge_pe                (merge_data_o_1_19),
    .ready_i_merge_pe               (merge_ready_i_1_19),

    .valid_i_gather_pe              (gather_valid_i_1_19),
    .data_i_gather_pe               (gather_data_i_1_19),
    .ready_o_gather_pe              (gather_ready_o_1_19),
    .valid_o_gather_pe              (gather_valid_o_1_19),
    .data_o_gather_pe               (gather_data_o_1_19),
    .ready_i_gather_pe              (gather_ready_i_1_19),

    .credit_upd                     (credit_upd[1][19])
);


network_interface #(
    .cast_out                       (cast_out_1_20),
    .gather_out                     (gather_out_1_20),
    .cast_sid                       (cast_sid_1_20),
    .gather_sid                     (gather_sid_1_20)
)ni_1_20(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[1][20]),
    .data_i_cast_nw                 (data_o_cast_nw[1][20]),
    .ready_o_cast_nw                (ready_i_cast_nw[1][20]),
    .valid_o_cast_nw                (valid_i_cast_nw[1][20]),
    .data_o_cast_nw                 (data_i_cast_nw[1][20]),
    .ready_i_cast_nw                (ready_o_cast_nw[1][20]),

    .valid_i_gather_nw              (valid_o_gather_nw[1][20]),
    .data_i_gather_nw               (data_o_gather_nw[1][20]),
    .ready_o_gather_nw              (ready_i_gather_nw[1][20]),
    .valid_o_gather_nw              (valid_i_gather_nw[1][20]),
    .data_o_gather_nw               (data_i_gather_nw[1][20]),
    .ready_i_gather_nw              (ready_o_gather_nw[1][20]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[1][20]),
    .data_i_merge_nw                (data_o_merge_nw[1][20]),
    .ready_o_merge_nw               (ready_i_merge_nw[1][20]),
    .valid_o_merge_nw               (valid_i_merge_nw[1][20]),
    .data_o_merge_nw                (data_i_merge_nw[1][20]),
    .ready_i_merge_nw               (ready_o_merge_nw[1][20]),

    .valid_i_cast_pe                (cast_valid_i_1_20),
    .data_i_cast_pe                 (cast_data_i_1_20),
    .ready_o_cast_pe                (cast_ready_o_1_20),
    .valid_o_cast_pe                (cast_valid_o_1_20),
    .data_o_cast_pe                 (cast_data_o_1_20),
    .ready_i_cast_pe                (cast_ready_i_1_20),

    .valid_i_merge_pe               (merge_valid_i_1_20),
    .data_i_merge_pe                (merge_data_i_1_20),
    .ready_o_merge_pe               (merge_ready_o_1_20),
    .valid_o_merge_pe               (merge_valid_o_1_20),
    .data_o_merge_pe                (merge_data_o_1_20),
    .ready_i_merge_pe               (merge_ready_i_1_20),

    .valid_i_gather_pe              (gather_valid_i_1_20),
    .data_i_gather_pe               (gather_data_i_1_20),
    .ready_o_gather_pe              (gather_ready_o_1_20),
    .valid_o_gather_pe              (gather_valid_o_1_20),
    .data_o_gather_pe               (gather_data_o_1_20),
    .ready_i_gather_pe              (gather_ready_i_1_20),

    .credit_upd                     (credit_upd[1][20])
);


network_interface #(
    .cast_out                       (cast_out_1_21),
    .gather_out                     (gather_out_1_21),
    .cast_sid                       (cast_sid_1_21),
    .gather_sid                     (gather_sid_1_21)
)ni_1_21(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[1][21]),
    .data_i_cast_nw                 (data_o_cast_nw[1][21]),
    .ready_o_cast_nw                (ready_i_cast_nw[1][21]),
    .valid_o_cast_nw                (valid_i_cast_nw[1][21]),
    .data_o_cast_nw                 (data_i_cast_nw[1][21]),
    .ready_i_cast_nw                (ready_o_cast_nw[1][21]),

    .valid_i_gather_nw              (valid_o_gather_nw[1][21]),
    .data_i_gather_nw               (data_o_gather_nw[1][21]),
    .ready_o_gather_nw              (ready_i_gather_nw[1][21]),
    .valid_o_gather_nw              (valid_i_gather_nw[1][21]),
    .data_o_gather_nw               (data_i_gather_nw[1][21]),
    .ready_i_gather_nw              (ready_o_gather_nw[1][21]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[1][21]),
    .data_i_merge_nw                (data_o_merge_nw[1][21]),
    .ready_o_merge_nw               (ready_i_merge_nw[1][21]),
    .valid_o_merge_nw               (valid_i_merge_nw[1][21]),
    .data_o_merge_nw                (data_i_merge_nw[1][21]),
    .ready_i_merge_nw               (ready_o_merge_nw[1][21]),

    .valid_i_cast_pe                (cast_valid_i_1_21),
    .data_i_cast_pe                 (cast_data_i_1_21),
    .ready_o_cast_pe                (cast_ready_o_1_21),
    .valid_o_cast_pe                (cast_valid_o_1_21),
    .data_o_cast_pe                 (cast_data_o_1_21),
    .ready_i_cast_pe                (cast_ready_i_1_21),

    .valid_i_merge_pe               (merge_valid_i_1_21),
    .data_i_merge_pe                (merge_data_i_1_21),
    .ready_o_merge_pe               (merge_ready_o_1_21),
    .valid_o_merge_pe               (merge_valid_o_1_21),
    .data_o_merge_pe                (merge_data_o_1_21),
    .ready_i_merge_pe               (merge_ready_i_1_21),

    .valid_i_gather_pe              (gather_valid_i_1_21),
    .data_i_gather_pe               (gather_data_i_1_21),
    .ready_o_gather_pe              (gather_ready_o_1_21),
    .valid_o_gather_pe              (gather_valid_o_1_21),
    .data_o_gather_pe               (gather_data_o_1_21),
    .ready_i_gather_pe              (gather_ready_i_1_21),

    .credit_upd                     (credit_upd[1][21])
);


network_interface #(
    .cast_out                       (cast_out_1_22),
    .gather_out                     (gather_out_1_22),
    .cast_sid                       (cast_sid_1_22),
    .gather_sid                     (gather_sid_1_22)
)ni_1_22(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[1][22]),
    .data_i_cast_nw                 (data_o_cast_nw[1][22]),
    .ready_o_cast_nw                (ready_i_cast_nw[1][22]),
    .valid_o_cast_nw                (valid_i_cast_nw[1][22]),
    .data_o_cast_nw                 (data_i_cast_nw[1][22]),
    .ready_i_cast_nw                (ready_o_cast_nw[1][22]),

    .valid_i_gather_nw              (valid_o_gather_nw[1][22]),
    .data_i_gather_nw               (data_o_gather_nw[1][22]),
    .ready_o_gather_nw              (ready_i_gather_nw[1][22]),
    .valid_o_gather_nw              (valid_i_gather_nw[1][22]),
    .data_o_gather_nw               (data_i_gather_nw[1][22]),
    .ready_i_gather_nw              (ready_o_gather_nw[1][22]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[1][22]),
    .data_i_merge_nw                (data_o_merge_nw[1][22]),
    .ready_o_merge_nw               (ready_i_merge_nw[1][22]),
    .valid_o_merge_nw               (valid_i_merge_nw[1][22]),
    .data_o_merge_nw                (data_i_merge_nw[1][22]),
    .ready_i_merge_nw               (ready_o_merge_nw[1][22]),

    .valid_i_cast_pe                (cast_valid_i_1_22),
    .data_i_cast_pe                 (cast_data_i_1_22),
    .ready_o_cast_pe                (cast_ready_o_1_22),
    .valid_o_cast_pe                (cast_valid_o_1_22),
    .data_o_cast_pe                 (cast_data_o_1_22),
    .ready_i_cast_pe                (cast_ready_i_1_22),

    .valid_i_merge_pe               (merge_valid_i_1_22),
    .data_i_merge_pe                (merge_data_i_1_22),
    .ready_o_merge_pe               (merge_ready_o_1_22),
    .valid_o_merge_pe               (merge_valid_o_1_22),
    .data_o_merge_pe                (merge_data_o_1_22),
    .ready_i_merge_pe               (merge_ready_i_1_22),

    .valid_i_gather_pe              (gather_valid_i_1_22),
    .data_i_gather_pe               (gather_data_i_1_22),
    .ready_o_gather_pe              (gather_ready_o_1_22),
    .valid_o_gather_pe              (gather_valid_o_1_22),
    .data_o_gather_pe               (gather_data_o_1_22),
    .ready_i_gather_pe              (gather_ready_i_1_22),

    .credit_upd                     (credit_upd[1][22])
);


network_interface #(
    .cast_out                       (cast_out_1_23),
    .gather_out                     (gather_out_1_23),
    .cast_sid                       (cast_sid_1_23),
    .gather_sid                     (gather_sid_1_23)
)ni_1_23(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[1][23]),
    .data_i_cast_nw                 (data_o_cast_nw[1][23]),
    .ready_o_cast_nw                (ready_i_cast_nw[1][23]),
    .valid_o_cast_nw                (valid_i_cast_nw[1][23]),
    .data_o_cast_nw                 (data_i_cast_nw[1][23]),
    .ready_i_cast_nw                (ready_o_cast_nw[1][23]),

    .valid_i_gather_nw              (valid_o_gather_nw[1][23]),
    .data_i_gather_nw               (data_o_gather_nw[1][23]),
    .ready_o_gather_nw              (ready_i_gather_nw[1][23]),
    .valid_o_gather_nw              (valid_i_gather_nw[1][23]),
    .data_o_gather_nw               (data_i_gather_nw[1][23]),
    .ready_i_gather_nw              (ready_o_gather_nw[1][23]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[1][23]),
    .data_i_merge_nw                (data_o_merge_nw[1][23]),
    .ready_o_merge_nw               (ready_i_merge_nw[1][23]),
    .valid_o_merge_nw               (valid_i_merge_nw[1][23]),
    .data_o_merge_nw                (data_i_merge_nw[1][23]),
    .ready_i_merge_nw               (ready_o_merge_nw[1][23]),

    .valid_i_cast_pe                (cast_valid_i_1_23),
    .data_i_cast_pe                 (cast_data_i_1_23),
    .ready_o_cast_pe                (cast_ready_o_1_23),
    .valid_o_cast_pe                (cast_valid_o_1_23),
    .data_o_cast_pe                 (cast_data_o_1_23),
    .ready_i_cast_pe                (cast_ready_i_1_23),

    .valid_i_merge_pe               (merge_valid_i_1_23),
    .data_i_merge_pe                (merge_data_i_1_23),
    .ready_o_merge_pe               (merge_ready_o_1_23),
    .valid_o_merge_pe               (merge_valid_o_1_23),
    .data_o_merge_pe                (merge_data_o_1_23),
    .ready_i_merge_pe               (merge_ready_i_1_23),

    .valid_i_gather_pe              (gather_valid_i_1_23),
    .data_i_gather_pe               (gather_data_i_1_23),
    .ready_o_gather_pe              (gather_ready_o_1_23),
    .valid_o_gather_pe              (gather_valid_o_1_23),
    .data_o_gather_pe               (gather_data_o_1_23),
    .ready_i_gather_pe              (gather_ready_i_1_23),

    .credit_upd                     (credit_upd[1][23])
);


network_interface #(
    .cast_out                       (cast_out_1_24),
    .gather_out                     (gather_out_1_24),
    .cast_sid                       (cast_sid_1_24),
    .gather_sid                     (gather_sid_1_24)
)ni_1_24(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[1][24]),
    .data_i_cast_nw                 (data_o_cast_nw[1][24]),
    .ready_o_cast_nw                (ready_i_cast_nw[1][24]),
    .valid_o_cast_nw                (valid_i_cast_nw[1][24]),
    .data_o_cast_nw                 (data_i_cast_nw[1][24]),
    .ready_i_cast_nw                (ready_o_cast_nw[1][24]),

    .valid_i_gather_nw              (valid_o_gather_nw[1][24]),
    .data_i_gather_nw               (data_o_gather_nw[1][24]),
    .ready_o_gather_nw              (ready_i_gather_nw[1][24]),
    .valid_o_gather_nw              (valid_i_gather_nw[1][24]),
    .data_o_gather_nw               (data_i_gather_nw[1][24]),
    .ready_i_gather_nw              (ready_o_gather_nw[1][24]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[1][24]),
    .data_i_merge_nw                (data_o_merge_nw[1][24]),
    .ready_o_merge_nw               (ready_i_merge_nw[1][24]),
    .valid_o_merge_nw               (valid_i_merge_nw[1][24]),
    .data_o_merge_nw                (data_i_merge_nw[1][24]),
    .ready_i_merge_nw               (ready_o_merge_nw[1][24]),

    .valid_i_cast_pe                (cast_valid_i_1_24),
    .data_i_cast_pe                 (cast_data_i_1_24),
    .ready_o_cast_pe                (cast_ready_o_1_24),
    .valid_o_cast_pe                (cast_valid_o_1_24),
    .data_o_cast_pe                 (cast_data_o_1_24),
    .ready_i_cast_pe                (cast_ready_i_1_24),

    .valid_i_merge_pe               (merge_valid_i_1_24),
    .data_i_merge_pe                (merge_data_i_1_24),
    .ready_o_merge_pe               (merge_ready_o_1_24),
    .valid_o_merge_pe               (merge_valid_o_1_24),
    .data_o_merge_pe                (merge_data_o_1_24),
    .ready_i_merge_pe               (merge_ready_i_1_24),

    .valid_i_gather_pe              (gather_valid_i_1_24),
    .data_i_gather_pe               (gather_data_i_1_24),
    .ready_o_gather_pe              (gather_ready_o_1_24),
    .valid_o_gather_pe              (gather_valid_o_1_24),
    .data_o_gather_pe               (gather_data_o_1_24),
    .ready_i_gather_pe              (gather_ready_i_1_24),

    .credit_upd                     (credit_upd[1][24])
);


network_interface #(
    .cast_out                       (cast_out_2_0),
    .gather_out                     (gather_out_2_0),
    .cast_sid                       (cast_sid_2_0),
    .gather_sid                     (gather_sid_2_0)
)ni_2_0(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[2][0]),
    .data_i_cast_nw                 (data_o_cast_nw[2][0]),
    .ready_o_cast_nw                (ready_i_cast_nw[2][0]),
    .valid_o_cast_nw                (valid_i_cast_nw[2][0]),
    .data_o_cast_nw                 (data_i_cast_nw[2][0]),
    .ready_i_cast_nw                (ready_o_cast_nw[2][0]),

    .valid_i_gather_nw              (valid_o_gather_nw[2][0]),
    .data_i_gather_nw               (data_o_gather_nw[2][0]),
    .ready_o_gather_nw              (ready_i_gather_nw[2][0]),
    .valid_o_gather_nw              (valid_i_gather_nw[2][0]),
    .data_o_gather_nw               (data_i_gather_nw[2][0]),
    .ready_i_gather_nw              (ready_o_gather_nw[2][0]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[2][0]),
    .data_i_merge_nw                (data_o_merge_nw[2][0]),
    .ready_o_merge_nw               (ready_i_merge_nw[2][0]),
    .valid_o_merge_nw               (valid_i_merge_nw[2][0]),
    .data_o_merge_nw                (data_i_merge_nw[2][0]),
    .ready_i_merge_nw               (ready_o_merge_nw[2][0]),

    .valid_i_cast_pe                (cast_valid_i_2_0),
    .data_i_cast_pe                 (cast_data_i_2_0),
    .ready_o_cast_pe                (cast_ready_o_2_0),
    .valid_o_cast_pe                (cast_valid_o_2_0),
    .data_o_cast_pe                 (cast_data_o_2_0),
    .ready_i_cast_pe                (cast_ready_i_2_0),

    .valid_i_merge_pe               (merge_valid_i_2_0),
    .data_i_merge_pe                (merge_data_i_2_0),
    .ready_o_merge_pe               (merge_ready_o_2_0),
    .valid_o_merge_pe               (merge_valid_o_2_0),
    .data_o_merge_pe                (merge_data_o_2_0),
    .ready_i_merge_pe               (merge_ready_i_2_0),

    .valid_i_gather_pe              (gather_valid_i_2_0),
    .data_i_gather_pe               (gather_data_i_2_0),
    .ready_o_gather_pe              (gather_ready_o_2_0),
    .valid_o_gather_pe              (gather_valid_o_2_0),
    .data_o_gather_pe               (gather_data_o_2_0),
    .ready_i_gather_pe              (gather_ready_i_2_0),

    .credit_upd                     (credit_upd[2][0])
);


network_interface #(
    .cast_out                       (cast_out_2_1),
    .gather_out                     (gather_out_2_1),
    .cast_sid                       (cast_sid_2_1),
    .gather_sid                     (gather_sid_2_1)
)ni_2_1(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[2][1]),
    .data_i_cast_nw                 (data_o_cast_nw[2][1]),
    .ready_o_cast_nw                (ready_i_cast_nw[2][1]),
    .valid_o_cast_nw                (valid_i_cast_nw[2][1]),
    .data_o_cast_nw                 (data_i_cast_nw[2][1]),
    .ready_i_cast_nw                (ready_o_cast_nw[2][1]),

    .valid_i_gather_nw              (valid_o_gather_nw[2][1]),
    .data_i_gather_nw               (data_o_gather_nw[2][1]),
    .ready_o_gather_nw              (ready_i_gather_nw[2][1]),
    .valid_o_gather_nw              (valid_i_gather_nw[2][1]),
    .data_o_gather_nw               (data_i_gather_nw[2][1]),
    .ready_i_gather_nw              (ready_o_gather_nw[2][1]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[2][1]),
    .data_i_merge_nw                (data_o_merge_nw[2][1]),
    .ready_o_merge_nw               (ready_i_merge_nw[2][1]),
    .valid_o_merge_nw               (valid_i_merge_nw[2][1]),
    .data_o_merge_nw                (data_i_merge_nw[2][1]),
    .ready_i_merge_nw               (ready_o_merge_nw[2][1]),

    .valid_i_cast_pe                (cast_valid_i_2_1),
    .data_i_cast_pe                 (cast_data_i_2_1),
    .ready_o_cast_pe                (cast_ready_o_2_1),
    .valid_o_cast_pe                (cast_valid_o_2_1),
    .data_o_cast_pe                 (cast_data_o_2_1),
    .ready_i_cast_pe                (cast_ready_i_2_1),

    .valid_i_merge_pe               (merge_valid_i_2_1),
    .data_i_merge_pe                (merge_data_i_2_1),
    .ready_o_merge_pe               (merge_ready_o_2_1),
    .valid_o_merge_pe               (merge_valid_o_2_1),
    .data_o_merge_pe                (merge_data_o_2_1),
    .ready_i_merge_pe               (merge_ready_i_2_1),

    .valid_i_gather_pe              (gather_valid_i_2_1),
    .data_i_gather_pe               (gather_data_i_2_1),
    .ready_o_gather_pe              (gather_ready_o_2_1),
    .valid_o_gather_pe              (gather_valid_o_2_1),
    .data_o_gather_pe               (gather_data_o_2_1),
    .ready_i_gather_pe              (gather_ready_i_2_1),

    .credit_upd                     (credit_upd[2][1])
);


network_interface #(
    .cast_out                       (cast_out_2_2),
    .gather_out                     (gather_out_2_2),
    .cast_sid                       (cast_sid_2_2),
    .gather_sid                     (gather_sid_2_2)
)ni_2_2(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[2][2]),
    .data_i_cast_nw                 (data_o_cast_nw[2][2]),
    .ready_o_cast_nw                (ready_i_cast_nw[2][2]),
    .valid_o_cast_nw                (valid_i_cast_nw[2][2]),
    .data_o_cast_nw                 (data_i_cast_nw[2][2]),
    .ready_i_cast_nw                (ready_o_cast_nw[2][2]),

    .valid_i_gather_nw              (valid_o_gather_nw[2][2]),
    .data_i_gather_nw               (data_o_gather_nw[2][2]),
    .ready_o_gather_nw              (ready_i_gather_nw[2][2]),
    .valid_o_gather_nw              (valid_i_gather_nw[2][2]),
    .data_o_gather_nw               (data_i_gather_nw[2][2]),
    .ready_i_gather_nw              (ready_o_gather_nw[2][2]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[2][2]),
    .data_i_merge_nw                (data_o_merge_nw[2][2]),
    .ready_o_merge_nw               (ready_i_merge_nw[2][2]),
    .valid_o_merge_nw               (valid_i_merge_nw[2][2]),
    .data_o_merge_nw                (data_i_merge_nw[2][2]),
    .ready_i_merge_nw               (ready_o_merge_nw[2][2]),

    .valid_i_cast_pe                (cast_valid_i_2_2),
    .data_i_cast_pe                 (cast_data_i_2_2),
    .ready_o_cast_pe                (cast_ready_o_2_2),
    .valid_o_cast_pe                (cast_valid_o_2_2),
    .data_o_cast_pe                 (cast_data_o_2_2),
    .ready_i_cast_pe                (cast_ready_i_2_2),

    .valid_i_merge_pe               (merge_valid_i_2_2),
    .data_i_merge_pe                (merge_data_i_2_2),
    .ready_o_merge_pe               (merge_ready_o_2_2),
    .valid_o_merge_pe               (merge_valid_o_2_2),
    .data_o_merge_pe                (merge_data_o_2_2),
    .ready_i_merge_pe               (merge_ready_i_2_2),

    .valid_i_gather_pe              (gather_valid_i_2_2),
    .data_i_gather_pe               (gather_data_i_2_2),
    .ready_o_gather_pe              (gather_ready_o_2_2),
    .valid_o_gather_pe              (gather_valid_o_2_2),
    .data_o_gather_pe               (gather_data_o_2_2),
    .ready_i_gather_pe              (gather_ready_i_2_2),

    .credit_upd                     (credit_upd[2][2])
);


network_interface #(
    .cast_out                       (cast_out_2_3),
    .gather_out                     (gather_out_2_3),
    .cast_sid                       (cast_sid_2_3),
    .gather_sid                     (gather_sid_2_3)
)ni_2_3(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[2][3]),
    .data_i_cast_nw                 (data_o_cast_nw[2][3]),
    .ready_o_cast_nw                (ready_i_cast_nw[2][3]),
    .valid_o_cast_nw                (valid_i_cast_nw[2][3]),
    .data_o_cast_nw                 (data_i_cast_nw[2][3]),
    .ready_i_cast_nw                (ready_o_cast_nw[2][3]),

    .valid_i_gather_nw              (valid_o_gather_nw[2][3]),
    .data_i_gather_nw               (data_o_gather_nw[2][3]),
    .ready_o_gather_nw              (ready_i_gather_nw[2][3]),
    .valid_o_gather_nw              (valid_i_gather_nw[2][3]),
    .data_o_gather_nw               (data_i_gather_nw[2][3]),
    .ready_i_gather_nw              (ready_o_gather_nw[2][3]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[2][3]),
    .data_i_merge_nw                (data_o_merge_nw[2][3]),
    .ready_o_merge_nw               (ready_i_merge_nw[2][3]),
    .valid_o_merge_nw               (valid_i_merge_nw[2][3]),
    .data_o_merge_nw                (data_i_merge_nw[2][3]),
    .ready_i_merge_nw               (ready_o_merge_nw[2][3]),

    .valid_i_cast_pe                (cast_valid_i_2_3),
    .data_i_cast_pe                 (cast_data_i_2_3),
    .ready_o_cast_pe                (cast_ready_o_2_3),
    .valid_o_cast_pe                (cast_valid_o_2_3),
    .data_o_cast_pe                 (cast_data_o_2_3),
    .ready_i_cast_pe                (cast_ready_i_2_3),

    .valid_i_merge_pe               (merge_valid_i_2_3),
    .data_i_merge_pe                (merge_data_i_2_3),
    .ready_o_merge_pe               (merge_ready_o_2_3),
    .valid_o_merge_pe               (merge_valid_o_2_3),
    .data_o_merge_pe                (merge_data_o_2_3),
    .ready_i_merge_pe               (merge_ready_i_2_3),

    .valid_i_gather_pe              (gather_valid_i_2_3),
    .data_i_gather_pe               (gather_data_i_2_3),
    .ready_o_gather_pe              (gather_ready_o_2_3),
    .valid_o_gather_pe              (gather_valid_o_2_3),
    .data_o_gather_pe               (gather_data_o_2_3),
    .ready_i_gather_pe              (gather_ready_i_2_3),

    .credit_upd                     (credit_upd[2][3])
);


network_interface #(
    .cast_out                       (cast_out_2_4),
    .gather_out                     (gather_out_2_4),
    .cast_sid                       (cast_sid_2_4),
    .gather_sid                     (gather_sid_2_4)
)ni_2_4(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[2][4]),
    .data_i_cast_nw                 (data_o_cast_nw[2][4]),
    .ready_o_cast_nw                (ready_i_cast_nw[2][4]),
    .valid_o_cast_nw                (valid_i_cast_nw[2][4]),
    .data_o_cast_nw                 (data_i_cast_nw[2][4]),
    .ready_i_cast_nw                (ready_o_cast_nw[2][4]),

    .valid_i_gather_nw              (valid_o_gather_nw[2][4]),
    .data_i_gather_nw               (data_o_gather_nw[2][4]),
    .ready_o_gather_nw              (ready_i_gather_nw[2][4]),
    .valid_o_gather_nw              (valid_i_gather_nw[2][4]),
    .data_o_gather_nw               (data_i_gather_nw[2][4]),
    .ready_i_gather_nw              (ready_o_gather_nw[2][4]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[2][4]),
    .data_i_merge_nw                (data_o_merge_nw[2][4]),
    .ready_o_merge_nw               (ready_i_merge_nw[2][4]),
    .valid_o_merge_nw               (valid_i_merge_nw[2][4]),
    .data_o_merge_nw                (data_i_merge_nw[2][4]),
    .ready_i_merge_nw               (ready_o_merge_nw[2][4]),

    .valid_i_cast_pe                (cast_valid_i_2_4),
    .data_i_cast_pe                 (cast_data_i_2_4),
    .ready_o_cast_pe                (cast_ready_o_2_4),
    .valid_o_cast_pe                (cast_valid_o_2_4),
    .data_o_cast_pe                 (cast_data_o_2_4),
    .ready_i_cast_pe                (cast_ready_i_2_4),

    .valid_i_merge_pe               (merge_valid_i_2_4),
    .data_i_merge_pe                (merge_data_i_2_4),
    .ready_o_merge_pe               (merge_ready_o_2_4),
    .valid_o_merge_pe               (merge_valid_o_2_4),
    .data_o_merge_pe                (merge_data_o_2_4),
    .ready_i_merge_pe               (merge_ready_i_2_4),

    .valid_i_gather_pe              (gather_valid_i_2_4),
    .data_i_gather_pe               (gather_data_i_2_4),
    .ready_o_gather_pe              (gather_ready_o_2_4),
    .valid_o_gather_pe              (gather_valid_o_2_4),
    .data_o_gather_pe               (gather_data_o_2_4),
    .ready_i_gather_pe              (gather_ready_i_2_4),

    .credit_upd                     (credit_upd[2][4])
);


network_interface #(
    .cast_out                       (cast_out_2_5),
    .gather_out                     (gather_out_2_5),
    .cast_sid                       (cast_sid_2_5),
    .gather_sid                     (gather_sid_2_5)
)ni_2_5(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[2][5]),
    .data_i_cast_nw                 (data_o_cast_nw[2][5]),
    .ready_o_cast_nw                (ready_i_cast_nw[2][5]),
    .valid_o_cast_nw                (valid_i_cast_nw[2][5]),
    .data_o_cast_nw                 (data_i_cast_nw[2][5]),
    .ready_i_cast_nw                (ready_o_cast_nw[2][5]),

    .valid_i_gather_nw              (valid_o_gather_nw[2][5]),
    .data_i_gather_nw               (data_o_gather_nw[2][5]),
    .ready_o_gather_nw              (ready_i_gather_nw[2][5]),
    .valid_o_gather_nw              (valid_i_gather_nw[2][5]),
    .data_o_gather_nw               (data_i_gather_nw[2][5]),
    .ready_i_gather_nw              (ready_o_gather_nw[2][5]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[2][5]),
    .data_i_merge_nw                (data_o_merge_nw[2][5]),
    .ready_o_merge_nw               (ready_i_merge_nw[2][5]),
    .valid_o_merge_nw               (valid_i_merge_nw[2][5]),
    .data_o_merge_nw                (data_i_merge_nw[2][5]),
    .ready_i_merge_nw               (ready_o_merge_nw[2][5]),

    .valid_i_cast_pe                (cast_valid_i_2_5),
    .data_i_cast_pe                 (cast_data_i_2_5),
    .ready_o_cast_pe                (cast_ready_o_2_5),
    .valid_o_cast_pe                (cast_valid_o_2_5),
    .data_o_cast_pe                 (cast_data_o_2_5),
    .ready_i_cast_pe                (cast_ready_i_2_5),

    .valid_i_merge_pe               (merge_valid_i_2_5),
    .data_i_merge_pe                (merge_data_i_2_5),
    .ready_o_merge_pe               (merge_ready_o_2_5),
    .valid_o_merge_pe               (merge_valid_o_2_5),
    .data_o_merge_pe                (merge_data_o_2_5),
    .ready_i_merge_pe               (merge_ready_i_2_5),

    .valid_i_gather_pe              (gather_valid_i_2_5),
    .data_i_gather_pe               (gather_data_i_2_5),
    .ready_o_gather_pe              (gather_ready_o_2_5),
    .valid_o_gather_pe              (gather_valid_o_2_5),
    .data_o_gather_pe               (gather_data_o_2_5),
    .ready_i_gather_pe              (gather_ready_i_2_5),

    .credit_upd                     (credit_upd[2][5])
);


network_interface #(
    .cast_out                       (cast_out_2_6),
    .gather_out                     (gather_out_2_6),
    .cast_sid                       (cast_sid_2_6),
    .gather_sid                     (gather_sid_2_6)
)ni_2_6(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[2][6]),
    .data_i_cast_nw                 (data_o_cast_nw[2][6]),
    .ready_o_cast_nw                (ready_i_cast_nw[2][6]),
    .valid_o_cast_nw                (valid_i_cast_nw[2][6]),
    .data_o_cast_nw                 (data_i_cast_nw[2][6]),
    .ready_i_cast_nw                (ready_o_cast_nw[2][6]),

    .valid_i_gather_nw              (valid_o_gather_nw[2][6]),
    .data_i_gather_nw               (data_o_gather_nw[2][6]),
    .ready_o_gather_nw              (ready_i_gather_nw[2][6]),
    .valid_o_gather_nw              (valid_i_gather_nw[2][6]),
    .data_o_gather_nw               (data_i_gather_nw[2][6]),
    .ready_i_gather_nw              (ready_o_gather_nw[2][6]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[2][6]),
    .data_i_merge_nw                (data_o_merge_nw[2][6]),
    .ready_o_merge_nw               (ready_i_merge_nw[2][6]),
    .valid_o_merge_nw               (valid_i_merge_nw[2][6]),
    .data_o_merge_nw                (data_i_merge_nw[2][6]),
    .ready_i_merge_nw               (ready_o_merge_nw[2][6]),

    .valid_i_cast_pe                (cast_valid_i_2_6),
    .data_i_cast_pe                 (cast_data_i_2_6),
    .ready_o_cast_pe                (cast_ready_o_2_6),
    .valid_o_cast_pe                (cast_valid_o_2_6),
    .data_o_cast_pe                 (cast_data_o_2_6),
    .ready_i_cast_pe                (cast_ready_i_2_6),

    .valid_i_merge_pe               (merge_valid_i_2_6),
    .data_i_merge_pe                (merge_data_i_2_6),
    .ready_o_merge_pe               (merge_ready_o_2_6),
    .valid_o_merge_pe               (merge_valid_o_2_6),
    .data_o_merge_pe                (merge_data_o_2_6),
    .ready_i_merge_pe               (merge_ready_i_2_6),

    .valid_i_gather_pe              (gather_valid_i_2_6),
    .data_i_gather_pe               (gather_data_i_2_6),
    .ready_o_gather_pe              (gather_ready_o_2_6),
    .valid_o_gather_pe              (gather_valid_o_2_6),
    .data_o_gather_pe               (gather_data_o_2_6),
    .ready_i_gather_pe              (gather_ready_i_2_6),

    .credit_upd                     (credit_upd[2][6])
);


network_interface #(
    .cast_out                       (cast_out_2_7),
    .gather_out                     (gather_out_2_7),
    .cast_sid                       (cast_sid_2_7),
    .gather_sid                     (gather_sid_2_7)
)ni_2_7(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[2][7]),
    .data_i_cast_nw                 (data_o_cast_nw[2][7]),
    .ready_o_cast_nw                (ready_i_cast_nw[2][7]),
    .valid_o_cast_nw                (valid_i_cast_nw[2][7]),
    .data_o_cast_nw                 (data_i_cast_nw[2][7]),
    .ready_i_cast_nw                (ready_o_cast_nw[2][7]),

    .valid_i_gather_nw              (valid_o_gather_nw[2][7]),
    .data_i_gather_nw               (data_o_gather_nw[2][7]),
    .ready_o_gather_nw              (ready_i_gather_nw[2][7]),
    .valid_o_gather_nw              (valid_i_gather_nw[2][7]),
    .data_o_gather_nw               (data_i_gather_nw[2][7]),
    .ready_i_gather_nw              (ready_o_gather_nw[2][7]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[2][7]),
    .data_i_merge_nw                (data_o_merge_nw[2][7]),
    .ready_o_merge_nw               (ready_i_merge_nw[2][7]),
    .valid_o_merge_nw               (valid_i_merge_nw[2][7]),
    .data_o_merge_nw                (data_i_merge_nw[2][7]),
    .ready_i_merge_nw               (ready_o_merge_nw[2][7]),

    .valid_i_cast_pe                (cast_valid_i_2_7),
    .data_i_cast_pe                 (cast_data_i_2_7),
    .ready_o_cast_pe                (cast_ready_o_2_7),
    .valid_o_cast_pe                (cast_valid_o_2_7),
    .data_o_cast_pe                 (cast_data_o_2_7),
    .ready_i_cast_pe                (cast_ready_i_2_7),

    .valid_i_merge_pe               (merge_valid_i_2_7),
    .data_i_merge_pe                (merge_data_i_2_7),
    .ready_o_merge_pe               (merge_ready_o_2_7),
    .valid_o_merge_pe               (merge_valid_o_2_7),
    .data_o_merge_pe                (merge_data_o_2_7),
    .ready_i_merge_pe               (merge_ready_i_2_7),

    .valid_i_gather_pe              (gather_valid_i_2_7),
    .data_i_gather_pe               (gather_data_i_2_7),
    .ready_o_gather_pe              (gather_ready_o_2_7),
    .valid_o_gather_pe              (gather_valid_o_2_7),
    .data_o_gather_pe               (gather_data_o_2_7),
    .ready_i_gather_pe              (gather_ready_i_2_7),

    .credit_upd                     (credit_upd[2][7])
);


network_interface #(
    .cast_out                       (cast_out_2_8),
    .gather_out                     (gather_out_2_8),
    .cast_sid                       (cast_sid_2_8),
    .gather_sid                     (gather_sid_2_8)
)ni_2_8(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[2][8]),
    .data_i_cast_nw                 (data_o_cast_nw[2][8]),
    .ready_o_cast_nw                (ready_i_cast_nw[2][8]),
    .valid_o_cast_nw                (valid_i_cast_nw[2][8]),
    .data_o_cast_nw                 (data_i_cast_nw[2][8]),
    .ready_i_cast_nw                (ready_o_cast_nw[2][8]),

    .valid_i_gather_nw              (valid_o_gather_nw[2][8]),
    .data_i_gather_nw               (data_o_gather_nw[2][8]),
    .ready_o_gather_nw              (ready_i_gather_nw[2][8]),
    .valid_o_gather_nw              (valid_i_gather_nw[2][8]),
    .data_o_gather_nw               (data_i_gather_nw[2][8]),
    .ready_i_gather_nw              (ready_o_gather_nw[2][8]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[2][8]),
    .data_i_merge_nw                (data_o_merge_nw[2][8]),
    .ready_o_merge_nw               (ready_i_merge_nw[2][8]),
    .valid_o_merge_nw               (valid_i_merge_nw[2][8]),
    .data_o_merge_nw                (data_i_merge_nw[2][8]),
    .ready_i_merge_nw               (ready_o_merge_nw[2][8]),

    .valid_i_cast_pe                (cast_valid_i_2_8),
    .data_i_cast_pe                 (cast_data_i_2_8),
    .ready_o_cast_pe                (cast_ready_o_2_8),
    .valid_o_cast_pe                (cast_valid_o_2_8),
    .data_o_cast_pe                 (cast_data_o_2_8),
    .ready_i_cast_pe                (cast_ready_i_2_8),

    .valid_i_merge_pe               (merge_valid_i_2_8),
    .data_i_merge_pe                (merge_data_i_2_8),
    .ready_o_merge_pe               (merge_ready_o_2_8),
    .valid_o_merge_pe               (merge_valid_o_2_8),
    .data_o_merge_pe                (merge_data_o_2_8),
    .ready_i_merge_pe               (merge_ready_i_2_8),

    .valid_i_gather_pe              (gather_valid_i_2_8),
    .data_i_gather_pe               (gather_data_i_2_8),
    .ready_o_gather_pe              (gather_ready_o_2_8),
    .valid_o_gather_pe              (gather_valid_o_2_8),
    .data_o_gather_pe               (gather_data_o_2_8),
    .ready_i_gather_pe              (gather_ready_i_2_8),

    .credit_upd                     (credit_upd[2][8])
);


network_interface #(
    .cast_out                       (cast_out_2_9),
    .gather_out                     (gather_out_2_9),
    .cast_sid                       (cast_sid_2_9),
    .gather_sid                     (gather_sid_2_9)
)ni_2_9(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[2][9]),
    .data_i_cast_nw                 (data_o_cast_nw[2][9]),
    .ready_o_cast_nw                (ready_i_cast_nw[2][9]),
    .valid_o_cast_nw                (valid_i_cast_nw[2][9]),
    .data_o_cast_nw                 (data_i_cast_nw[2][9]),
    .ready_i_cast_nw                (ready_o_cast_nw[2][9]),

    .valid_i_gather_nw              (valid_o_gather_nw[2][9]),
    .data_i_gather_nw               (data_o_gather_nw[2][9]),
    .ready_o_gather_nw              (ready_i_gather_nw[2][9]),
    .valid_o_gather_nw              (valid_i_gather_nw[2][9]),
    .data_o_gather_nw               (data_i_gather_nw[2][9]),
    .ready_i_gather_nw              (ready_o_gather_nw[2][9]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[2][9]),
    .data_i_merge_nw                (data_o_merge_nw[2][9]),
    .ready_o_merge_nw               (ready_i_merge_nw[2][9]),
    .valid_o_merge_nw               (valid_i_merge_nw[2][9]),
    .data_o_merge_nw                (data_i_merge_nw[2][9]),
    .ready_i_merge_nw               (ready_o_merge_nw[2][9]),

    .valid_i_cast_pe                (cast_valid_i_2_9),
    .data_i_cast_pe                 (cast_data_i_2_9),
    .ready_o_cast_pe                (cast_ready_o_2_9),
    .valid_o_cast_pe                (cast_valid_o_2_9),
    .data_o_cast_pe                 (cast_data_o_2_9),
    .ready_i_cast_pe                (cast_ready_i_2_9),

    .valid_i_merge_pe               (merge_valid_i_2_9),
    .data_i_merge_pe                (merge_data_i_2_9),
    .ready_o_merge_pe               (merge_ready_o_2_9),
    .valid_o_merge_pe               (merge_valid_o_2_9),
    .data_o_merge_pe                (merge_data_o_2_9),
    .ready_i_merge_pe               (merge_ready_i_2_9),

    .valid_i_gather_pe              (gather_valid_i_2_9),
    .data_i_gather_pe               (gather_data_i_2_9),
    .ready_o_gather_pe              (gather_ready_o_2_9),
    .valid_o_gather_pe              (gather_valid_o_2_9),
    .data_o_gather_pe               (gather_data_o_2_9),
    .ready_i_gather_pe              (gather_ready_i_2_9),

    .credit_upd                     (credit_upd[2][9])
);


network_interface #(
    .cast_out                       (cast_out_2_10),
    .gather_out                     (gather_out_2_10),
    .cast_sid                       (cast_sid_2_10),
    .gather_sid                     (gather_sid_2_10)
)ni_2_10(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[2][10]),
    .data_i_cast_nw                 (data_o_cast_nw[2][10]),
    .ready_o_cast_nw                (ready_i_cast_nw[2][10]),
    .valid_o_cast_nw                (valid_i_cast_nw[2][10]),
    .data_o_cast_nw                 (data_i_cast_nw[2][10]),
    .ready_i_cast_nw                (ready_o_cast_nw[2][10]),

    .valid_i_gather_nw              (valid_o_gather_nw[2][10]),
    .data_i_gather_nw               (data_o_gather_nw[2][10]),
    .ready_o_gather_nw              (ready_i_gather_nw[2][10]),
    .valid_o_gather_nw              (valid_i_gather_nw[2][10]),
    .data_o_gather_nw               (data_i_gather_nw[2][10]),
    .ready_i_gather_nw              (ready_o_gather_nw[2][10]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[2][10]),
    .data_i_merge_nw                (data_o_merge_nw[2][10]),
    .ready_o_merge_nw               (ready_i_merge_nw[2][10]),
    .valid_o_merge_nw               (valid_i_merge_nw[2][10]),
    .data_o_merge_nw                (data_i_merge_nw[2][10]),
    .ready_i_merge_nw               (ready_o_merge_nw[2][10]),

    .valid_i_cast_pe                (cast_valid_i_2_10),
    .data_i_cast_pe                 (cast_data_i_2_10),
    .ready_o_cast_pe                (cast_ready_o_2_10),
    .valid_o_cast_pe                (cast_valid_o_2_10),
    .data_o_cast_pe                 (cast_data_o_2_10),
    .ready_i_cast_pe                (cast_ready_i_2_10),

    .valid_i_merge_pe               (merge_valid_i_2_10),
    .data_i_merge_pe                (merge_data_i_2_10),
    .ready_o_merge_pe               (merge_ready_o_2_10),
    .valid_o_merge_pe               (merge_valid_o_2_10),
    .data_o_merge_pe                (merge_data_o_2_10),
    .ready_i_merge_pe               (merge_ready_i_2_10),

    .valid_i_gather_pe              (gather_valid_i_2_10),
    .data_i_gather_pe               (gather_data_i_2_10),
    .ready_o_gather_pe              (gather_ready_o_2_10),
    .valid_o_gather_pe              (gather_valid_o_2_10),
    .data_o_gather_pe               (gather_data_o_2_10),
    .ready_i_gather_pe              (gather_ready_i_2_10),

    .credit_upd                     (credit_upd[2][10])
);


network_interface #(
    .cast_out                       (cast_out_2_11),
    .gather_out                     (gather_out_2_11),
    .cast_sid                       (cast_sid_2_11),
    .gather_sid                     (gather_sid_2_11)
)ni_2_11(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[2][11]),
    .data_i_cast_nw                 (data_o_cast_nw[2][11]),
    .ready_o_cast_nw                (ready_i_cast_nw[2][11]),
    .valid_o_cast_nw                (valid_i_cast_nw[2][11]),
    .data_o_cast_nw                 (data_i_cast_nw[2][11]),
    .ready_i_cast_nw                (ready_o_cast_nw[2][11]),

    .valid_i_gather_nw              (valid_o_gather_nw[2][11]),
    .data_i_gather_nw               (data_o_gather_nw[2][11]),
    .ready_o_gather_nw              (ready_i_gather_nw[2][11]),
    .valid_o_gather_nw              (valid_i_gather_nw[2][11]),
    .data_o_gather_nw               (data_i_gather_nw[2][11]),
    .ready_i_gather_nw              (ready_o_gather_nw[2][11]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[2][11]),
    .data_i_merge_nw                (data_o_merge_nw[2][11]),
    .ready_o_merge_nw               (ready_i_merge_nw[2][11]),
    .valid_o_merge_nw               (valid_i_merge_nw[2][11]),
    .data_o_merge_nw                (data_i_merge_nw[2][11]),
    .ready_i_merge_nw               (ready_o_merge_nw[2][11]),

    .valid_i_cast_pe                (cast_valid_i_2_11),
    .data_i_cast_pe                 (cast_data_i_2_11),
    .ready_o_cast_pe                (cast_ready_o_2_11),
    .valid_o_cast_pe                (cast_valid_o_2_11),
    .data_o_cast_pe                 (cast_data_o_2_11),
    .ready_i_cast_pe                (cast_ready_i_2_11),

    .valid_i_merge_pe               (merge_valid_i_2_11),
    .data_i_merge_pe                (merge_data_i_2_11),
    .ready_o_merge_pe               (merge_ready_o_2_11),
    .valid_o_merge_pe               (merge_valid_o_2_11),
    .data_o_merge_pe                (merge_data_o_2_11),
    .ready_i_merge_pe               (merge_ready_i_2_11),

    .valid_i_gather_pe              (gather_valid_i_2_11),
    .data_i_gather_pe               (gather_data_i_2_11),
    .ready_o_gather_pe              (gather_ready_o_2_11),
    .valid_o_gather_pe              (gather_valid_o_2_11),
    .data_o_gather_pe               (gather_data_o_2_11),
    .ready_i_gather_pe              (gather_ready_i_2_11),

    .credit_upd                     (credit_upd[2][11])
);


network_interface #(
    .cast_out                       (cast_out_2_12),
    .gather_out                     (gather_out_2_12),
    .cast_sid                       (cast_sid_2_12),
    .gather_sid                     (gather_sid_2_12)
)ni_2_12(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[2][12]),
    .data_i_cast_nw                 (data_o_cast_nw[2][12]),
    .ready_o_cast_nw                (ready_i_cast_nw[2][12]),
    .valid_o_cast_nw                (valid_i_cast_nw[2][12]),
    .data_o_cast_nw                 (data_i_cast_nw[2][12]),
    .ready_i_cast_nw                (ready_o_cast_nw[2][12]),

    .valid_i_gather_nw              (valid_o_gather_nw[2][12]),
    .data_i_gather_nw               (data_o_gather_nw[2][12]),
    .ready_o_gather_nw              (ready_i_gather_nw[2][12]),
    .valid_o_gather_nw              (valid_i_gather_nw[2][12]),
    .data_o_gather_nw               (data_i_gather_nw[2][12]),
    .ready_i_gather_nw              (ready_o_gather_nw[2][12]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[2][12]),
    .data_i_merge_nw                (data_o_merge_nw[2][12]),
    .ready_o_merge_nw               (ready_i_merge_nw[2][12]),
    .valid_o_merge_nw               (valid_i_merge_nw[2][12]),
    .data_o_merge_nw                (data_i_merge_nw[2][12]),
    .ready_i_merge_nw               (ready_o_merge_nw[2][12]),

    .valid_i_cast_pe                (cast_valid_i_2_12),
    .data_i_cast_pe                 (cast_data_i_2_12),
    .ready_o_cast_pe                (cast_ready_o_2_12),
    .valid_o_cast_pe                (cast_valid_o_2_12),
    .data_o_cast_pe                 (cast_data_o_2_12),
    .ready_i_cast_pe                (cast_ready_i_2_12),

    .valid_i_merge_pe               (merge_valid_i_2_12),
    .data_i_merge_pe                (merge_data_i_2_12),
    .ready_o_merge_pe               (merge_ready_o_2_12),
    .valid_o_merge_pe               (merge_valid_o_2_12),
    .data_o_merge_pe                (merge_data_o_2_12),
    .ready_i_merge_pe               (merge_ready_i_2_12),

    .valid_i_gather_pe              (gather_valid_i_2_12),
    .data_i_gather_pe               (gather_data_i_2_12),
    .ready_o_gather_pe              (gather_ready_o_2_12),
    .valid_o_gather_pe              (gather_valid_o_2_12),
    .data_o_gather_pe               (gather_data_o_2_12),
    .ready_i_gather_pe              (gather_ready_i_2_12),

    .credit_upd                     (credit_upd[2][12])
);


network_interface #(
    .cast_out                       (cast_out_2_13),
    .gather_out                     (gather_out_2_13),
    .cast_sid                       (cast_sid_2_13),
    .gather_sid                     (gather_sid_2_13)
)ni_2_13(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[2][13]),
    .data_i_cast_nw                 (data_o_cast_nw[2][13]),
    .ready_o_cast_nw                (ready_i_cast_nw[2][13]),
    .valid_o_cast_nw                (valid_i_cast_nw[2][13]),
    .data_o_cast_nw                 (data_i_cast_nw[2][13]),
    .ready_i_cast_nw                (ready_o_cast_nw[2][13]),

    .valid_i_gather_nw              (valid_o_gather_nw[2][13]),
    .data_i_gather_nw               (data_o_gather_nw[2][13]),
    .ready_o_gather_nw              (ready_i_gather_nw[2][13]),
    .valid_o_gather_nw              (valid_i_gather_nw[2][13]),
    .data_o_gather_nw               (data_i_gather_nw[2][13]),
    .ready_i_gather_nw              (ready_o_gather_nw[2][13]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[2][13]),
    .data_i_merge_nw                (data_o_merge_nw[2][13]),
    .ready_o_merge_nw               (ready_i_merge_nw[2][13]),
    .valid_o_merge_nw               (valid_i_merge_nw[2][13]),
    .data_o_merge_nw                (data_i_merge_nw[2][13]),
    .ready_i_merge_nw               (ready_o_merge_nw[2][13]),

    .valid_i_cast_pe                (cast_valid_i_2_13),
    .data_i_cast_pe                 (cast_data_i_2_13),
    .ready_o_cast_pe                (cast_ready_o_2_13),
    .valid_o_cast_pe                (cast_valid_o_2_13),
    .data_o_cast_pe                 (cast_data_o_2_13),
    .ready_i_cast_pe                (cast_ready_i_2_13),

    .valid_i_merge_pe               (merge_valid_i_2_13),
    .data_i_merge_pe                (merge_data_i_2_13),
    .ready_o_merge_pe               (merge_ready_o_2_13),
    .valid_o_merge_pe               (merge_valid_o_2_13),
    .data_o_merge_pe                (merge_data_o_2_13),
    .ready_i_merge_pe               (merge_ready_i_2_13),

    .valid_i_gather_pe              (gather_valid_i_2_13),
    .data_i_gather_pe               (gather_data_i_2_13),
    .ready_o_gather_pe              (gather_ready_o_2_13),
    .valid_o_gather_pe              (gather_valid_o_2_13),
    .data_o_gather_pe               (gather_data_o_2_13),
    .ready_i_gather_pe              (gather_ready_i_2_13),

    .credit_upd                     (credit_upd[2][13])
);


network_interface #(
    .cast_out                       (cast_out_2_14),
    .gather_out                     (gather_out_2_14),
    .cast_sid                       (cast_sid_2_14),
    .gather_sid                     (gather_sid_2_14)
)ni_2_14(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[2][14]),
    .data_i_cast_nw                 (data_o_cast_nw[2][14]),
    .ready_o_cast_nw                (ready_i_cast_nw[2][14]),
    .valid_o_cast_nw                (valid_i_cast_nw[2][14]),
    .data_o_cast_nw                 (data_i_cast_nw[2][14]),
    .ready_i_cast_nw                (ready_o_cast_nw[2][14]),

    .valid_i_gather_nw              (valid_o_gather_nw[2][14]),
    .data_i_gather_nw               (data_o_gather_nw[2][14]),
    .ready_o_gather_nw              (ready_i_gather_nw[2][14]),
    .valid_o_gather_nw              (valid_i_gather_nw[2][14]),
    .data_o_gather_nw               (data_i_gather_nw[2][14]),
    .ready_i_gather_nw              (ready_o_gather_nw[2][14]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[2][14]),
    .data_i_merge_nw                (data_o_merge_nw[2][14]),
    .ready_o_merge_nw               (ready_i_merge_nw[2][14]),
    .valid_o_merge_nw               (valid_i_merge_nw[2][14]),
    .data_o_merge_nw                (data_i_merge_nw[2][14]),
    .ready_i_merge_nw               (ready_o_merge_nw[2][14]),

    .valid_i_cast_pe                (cast_valid_i_2_14),
    .data_i_cast_pe                 (cast_data_i_2_14),
    .ready_o_cast_pe                (cast_ready_o_2_14),
    .valid_o_cast_pe                (cast_valid_o_2_14),
    .data_o_cast_pe                 (cast_data_o_2_14),
    .ready_i_cast_pe                (cast_ready_i_2_14),

    .valid_i_merge_pe               (merge_valid_i_2_14),
    .data_i_merge_pe                (merge_data_i_2_14),
    .ready_o_merge_pe               (merge_ready_o_2_14),
    .valid_o_merge_pe               (merge_valid_o_2_14),
    .data_o_merge_pe                (merge_data_o_2_14),
    .ready_i_merge_pe               (merge_ready_i_2_14),

    .valid_i_gather_pe              (gather_valid_i_2_14),
    .data_i_gather_pe               (gather_data_i_2_14),
    .ready_o_gather_pe              (gather_ready_o_2_14),
    .valid_o_gather_pe              (gather_valid_o_2_14),
    .data_o_gather_pe               (gather_data_o_2_14),
    .ready_i_gather_pe              (gather_ready_i_2_14),

    .credit_upd                     (credit_upd[2][14])
);


network_interface #(
    .cast_out                       (cast_out_2_15),
    .gather_out                     (gather_out_2_15),
    .cast_sid                       (cast_sid_2_15),
    .gather_sid                     (gather_sid_2_15)
)ni_2_15(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[2][15]),
    .data_i_cast_nw                 (data_o_cast_nw[2][15]),
    .ready_o_cast_nw                (ready_i_cast_nw[2][15]),
    .valid_o_cast_nw                (valid_i_cast_nw[2][15]),
    .data_o_cast_nw                 (data_i_cast_nw[2][15]),
    .ready_i_cast_nw                (ready_o_cast_nw[2][15]),

    .valid_i_gather_nw              (valid_o_gather_nw[2][15]),
    .data_i_gather_nw               (data_o_gather_nw[2][15]),
    .ready_o_gather_nw              (ready_i_gather_nw[2][15]),
    .valid_o_gather_nw              (valid_i_gather_nw[2][15]),
    .data_o_gather_nw               (data_i_gather_nw[2][15]),
    .ready_i_gather_nw              (ready_o_gather_nw[2][15]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[2][15]),
    .data_i_merge_nw                (data_o_merge_nw[2][15]),
    .ready_o_merge_nw               (ready_i_merge_nw[2][15]),
    .valid_o_merge_nw               (valid_i_merge_nw[2][15]),
    .data_o_merge_nw                (data_i_merge_nw[2][15]),
    .ready_i_merge_nw               (ready_o_merge_nw[2][15]),

    .valid_i_cast_pe                (cast_valid_i_2_15),
    .data_i_cast_pe                 (cast_data_i_2_15),
    .ready_o_cast_pe                (cast_ready_o_2_15),
    .valid_o_cast_pe                (cast_valid_o_2_15),
    .data_o_cast_pe                 (cast_data_o_2_15),
    .ready_i_cast_pe                (cast_ready_i_2_15),

    .valid_i_merge_pe               (merge_valid_i_2_15),
    .data_i_merge_pe                (merge_data_i_2_15),
    .ready_o_merge_pe               (merge_ready_o_2_15),
    .valid_o_merge_pe               (merge_valid_o_2_15),
    .data_o_merge_pe                (merge_data_o_2_15),
    .ready_i_merge_pe               (merge_ready_i_2_15),

    .valid_i_gather_pe              (gather_valid_i_2_15),
    .data_i_gather_pe               (gather_data_i_2_15),
    .ready_o_gather_pe              (gather_ready_o_2_15),
    .valid_o_gather_pe              (gather_valid_o_2_15),
    .data_o_gather_pe               (gather_data_o_2_15),
    .ready_i_gather_pe              (gather_ready_i_2_15),

    .credit_upd                     (credit_upd[2][15])
);


network_interface #(
    .cast_out                       (cast_out_2_16),
    .gather_out                     (gather_out_2_16),
    .cast_sid                       (cast_sid_2_16),
    .gather_sid                     (gather_sid_2_16)
)ni_2_16(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[2][16]),
    .data_i_cast_nw                 (data_o_cast_nw[2][16]),
    .ready_o_cast_nw                (ready_i_cast_nw[2][16]),
    .valid_o_cast_nw                (valid_i_cast_nw[2][16]),
    .data_o_cast_nw                 (data_i_cast_nw[2][16]),
    .ready_i_cast_nw                (ready_o_cast_nw[2][16]),

    .valid_i_gather_nw              (valid_o_gather_nw[2][16]),
    .data_i_gather_nw               (data_o_gather_nw[2][16]),
    .ready_o_gather_nw              (ready_i_gather_nw[2][16]),
    .valid_o_gather_nw              (valid_i_gather_nw[2][16]),
    .data_o_gather_nw               (data_i_gather_nw[2][16]),
    .ready_i_gather_nw              (ready_o_gather_nw[2][16]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[2][16]),
    .data_i_merge_nw                (data_o_merge_nw[2][16]),
    .ready_o_merge_nw               (ready_i_merge_nw[2][16]),
    .valid_o_merge_nw               (valid_i_merge_nw[2][16]),
    .data_o_merge_nw                (data_i_merge_nw[2][16]),
    .ready_i_merge_nw               (ready_o_merge_nw[2][16]),

    .valid_i_cast_pe                (cast_valid_i_2_16),
    .data_i_cast_pe                 (cast_data_i_2_16),
    .ready_o_cast_pe                (cast_ready_o_2_16),
    .valid_o_cast_pe                (cast_valid_o_2_16),
    .data_o_cast_pe                 (cast_data_o_2_16),
    .ready_i_cast_pe                (cast_ready_i_2_16),

    .valid_i_merge_pe               (merge_valid_i_2_16),
    .data_i_merge_pe                (merge_data_i_2_16),
    .ready_o_merge_pe               (merge_ready_o_2_16),
    .valid_o_merge_pe               (merge_valid_o_2_16),
    .data_o_merge_pe                (merge_data_o_2_16),
    .ready_i_merge_pe               (merge_ready_i_2_16),

    .valid_i_gather_pe              (gather_valid_i_2_16),
    .data_i_gather_pe               (gather_data_i_2_16),
    .ready_o_gather_pe              (gather_ready_o_2_16),
    .valid_o_gather_pe              (gather_valid_o_2_16),
    .data_o_gather_pe               (gather_data_o_2_16),
    .ready_i_gather_pe              (gather_ready_i_2_16),

    .credit_upd                     (credit_upd[2][16])
);


network_interface #(
    .cast_out                       (cast_out_2_17),
    .gather_out                     (gather_out_2_17),
    .cast_sid                       (cast_sid_2_17),
    .gather_sid                     (gather_sid_2_17)
)ni_2_17(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[2][17]),
    .data_i_cast_nw                 (data_o_cast_nw[2][17]),
    .ready_o_cast_nw                (ready_i_cast_nw[2][17]),
    .valid_o_cast_nw                (valid_i_cast_nw[2][17]),
    .data_o_cast_nw                 (data_i_cast_nw[2][17]),
    .ready_i_cast_nw                (ready_o_cast_nw[2][17]),

    .valid_i_gather_nw              (valid_o_gather_nw[2][17]),
    .data_i_gather_nw               (data_o_gather_nw[2][17]),
    .ready_o_gather_nw              (ready_i_gather_nw[2][17]),
    .valid_o_gather_nw              (valid_i_gather_nw[2][17]),
    .data_o_gather_nw               (data_i_gather_nw[2][17]),
    .ready_i_gather_nw              (ready_o_gather_nw[2][17]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[2][17]),
    .data_i_merge_nw                (data_o_merge_nw[2][17]),
    .ready_o_merge_nw               (ready_i_merge_nw[2][17]),
    .valid_o_merge_nw               (valid_i_merge_nw[2][17]),
    .data_o_merge_nw                (data_i_merge_nw[2][17]),
    .ready_i_merge_nw               (ready_o_merge_nw[2][17]),

    .valid_i_cast_pe                (cast_valid_i_2_17),
    .data_i_cast_pe                 (cast_data_i_2_17),
    .ready_o_cast_pe                (cast_ready_o_2_17),
    .valid_o_cast_pe                (cast_valid_o_2_17),
    .data_o_cast_pe                 (cast_data_o_2_17),
    .ready_i_cast_pe                (cast_ready_i_2_17),

    .valid_i_merge_pe               (merge_valid_i_2_17),
    .data_i_merge_pe                (merge_data_i_2_17),
    .ready_o_merge_pe               (merge_ready_o_2_17),
    .valid_o_merge_pe               (merge_valid_o_2_17),
    .data_o_merge_pe                (merge_data_o_2_17),
    .ready_i_merge_pe               (merge_ready_i_2_17),

    .valid_i_gather_pe              (gather_valid_i_2_17),
    .data_i_gather_pe               (gather_data_i_2_17),
    .ready_o_gather_pe              (gather_ready_o_2_17),
    .valid_o_gather_pe              (gather_valid_o_2_17),
    .data_o_gather_pe               (gather_data_o_2_17),
    .ready_i_gather_pe              (gather_ready_i_2_17),

    .credit_upd                     (credit_upd[2][17])
);


network_interface #(
    .cast_out                       (cast_out_2_18),
    .gather_out                     (gather_out_2_18),
    .cast_sid                       (cast_sid_2_18),
    .gather_sid                     (gather_sid_2_18)
)ni_2_18(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[2][18]),
    .data_i_cast_nw                 (data_o_cast_nw[2][18]),
    .ready_o_cast_nw                (ready_i_cast_nw[2][18]),
    .valid_o_cast_nw                (valid_i_cast_nw[2][18]),
    .data_o_cast_nw                 (data_i_cast_nw[2][18]),
    .ready_i_cast_nw                (ready_o_cast_nw[2][18]),

    .valid_i_gather_nw              (valid_o_gather_nw[2][18]),
    .data_i_gather_nw               (data_o_gather_nw[2][18]),
    .ready_o_gather_nw              (ready_i_gather_nw[2][18]),
    .valid_o_gather_nw              (valid_i_gather_nw[2][18]),
    .data_o_gather_nw               (data_i_gather_nw[2][18]),
    .ready_i_gather_nw              (ready_o_gather_nw[2][18]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[2][18]),
    .data_i_merge_nw                (data_o_merge_nw[2][18]),
    .ready_o_merge_nw               (ready_i_merge_nw[2][18]),
    .valid_o_merge_nw               (valid_i_merge_nw[2][18]),
    .data_o_merge_nw                (data_i_merge_nw[2][18]),
    .ready_i_merge_nw               (ready_o_merge_nw[2][18]),

    .valid_i_cast_pe                (cast_valid_i_2_18),
    .data_i_cast_pe                 (cast_data_i_2_18),
    .ready_o_cast_pe                (cast_ready_o_2_18),
    .valid_o_cast_pe                (cast_valid_o_2_18),
    .data_o_cast_pe                 (cast_data_o_2_18),
    .ready_i_cast_pe                (cast_ready_i_2_18),

    .valid_i_merge_pe               (merge_valid_i_2_18),
    .data_i_merge_pe                (merge_data_i_2_18),
    .ready_o_merge_pe               (merge_ready_o_2_18),
    .valid_o_merge_pe               (merge_valid_o_2_18),
    .data_o_merge_pe                (merge_data_o_2_18),
    .ready_i_merge_pe               (merge_ready_i_2_18),

    .valid_i_gather_pe              (gather_valid_i_2_18),
    .data_i_gather_pe               (gather_data_i_2_18),
    .ready_o_gather_pe              (gather_ready_o_2_18),
    .valid_o_gather_pe              (gather_valid_o_2_18),
    .data_o_gather_pe               (gather_data_o_2_18),
    .ready_i_gather_pe              (gather_ready_i_2_18),

    .credit_upd                     (credit_upd[2][18])
);


network_interface #(
    .cast_out                       (cast_out_2_19),
    .gather_out                     (gather_out_2_19),
    .cast_sid                       (cast_sid_2_19),
    .gather_sid                     (gather_sid_2_19)
)ni_2_19(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[2][19]),
    .data_i_cast_nw                 (data_o_cast_nw[2][19]),
    .ready_o_cast_nw                (ready_i_cast_nw[2][19]),
    .valid_o_cast_nw                (valid_i_cast_nw[2][19]),
    .data_o_cast_nw                 (data_i_cast_nw[2][19]),
    .ready_i_cast_nw                (ready_o_cast_nw[2][19]),

    .valid_i_gather_nw              (valid_o_gather_nw[2][19]),
    .data_i_gather_nw               (data_o_gather_nw[2][19]),
    .ready_o_gather_nw              (ready_i_gather_nw[2][19]),
    .valid_o_gather_nw              (valid_i_gather_nw[2][19]),
    .data_o_gather_nw               (data_i_gather_nw[2][19]),
    .ready_i_gather_nw              (ready_o_gather_nw[2][19]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[2][19]),
    .data_i_merge_nw                (data_o_merge_nw[2][19]),
    .ready_o_merge_nw               (ready_i_merge_nw[2][19]),
    .valid_o_merge_nw               (valid_i_merge_nw[2][19]),
    .data_o_merge_nw                (data_i_merge_nw[2][19]),
    .ready_i_merge_nw               (ready_o_merge_nw[2][19]),

    .valid_i_cast_pe                (cast_valid_i_2_19),
    .data_i_cast_pe                 (cast_data_i_2_19),
    .ready_o_cast_pe                (cast_ready_o_2_19),
    .valid_o_cast_pe                (cast_valid_o_2_19),
    .data_o_cast_pe                 (cast_data_o_2_19),
    .ready_i_cast_pe                (cast_ready_i_2_19),

    .valid_i_merge_pe               (merge_valid_i_2_19),
    .data_i_merge_pe                (merge_data_i_2_19),
    .ready_o_merge_pe               (merge_ready_o_2_19),
    .valid_o_merge_pe               (merge_valid_o_2_19),
    .data_o_merge_pe                (merge_data_o_2_19),
    .ready_i_merge_pe               (merge_ready_i_2_19),

    .valid_i_gather_pe              (gather_valid_i_2_19),
    .data_i_gather_pe               (gather_data_i_2_19),
    .ready_o_gather_pe              (gather_ready_o_2_19),
    .valid_o_gather_pe              (gather_valid_o_2_19),
    .data_o_gather_pe               (gather_data_o_2_19),
    .ready_i_gather_pe              (gather_ready_i_2_19),

    .credit_upd                     (credit_upd[2][19])
);


network_interface #(
    .cast_out                       (cast_out_2_20),
    .gather_out                     (gather_out_2_20),
    .cast_sid                       (cast_sid_2_20),
    .gather_sid                     (gather_sid_2_20)
)ni_2_20(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[2][20]),
    .data_i_cast_nw                 (data_o_cast_nw[2][20]),
    .ready_o_cast_nw                (ready_i_cast_nw[2][20]),
    .valid_o_cast_nw                (valid_i_cast_nw[2][20]),
    .data_o_cast_nw                 (data_i_cast_nw[2][20]),
    .ready_i_cast_nw                (ready_o_cast_nw[2][20]),

    .valid_i_gather_nw              (valid_o_gather_nw[2][20]),
    .data_i_gather_nw               (data_o_gather_nw[2][20]),
    .ready_o_gather_nw              (ready_i_gather_nw[2][20]),
    .valid_o_gather_nw              (valid_i_gather_nw[2][20]),
    .data_o_gather_nw               (data_i_gather_nw[2][20]),
    .ready_i_gather_nw              (ready_o_gather_nw[2][20]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[2][20]),
    .data_i_merge_nw                (data_o_merge_nw[2][20]),
    .ready_o_merge_nw               (ready_i_merge_nw[2][20]),
    .valid_o_merge_nw               (valid_i_merge_nw[2][20]),
    .data_o_merge_nw                (data_i_merge_nw[2][20]),
    .ready_i_merge_nw               (ready_o_merge_nw[2][20]),

    .valid_i_cast_pe                (cast_valid_i_2_20),
    .data_i_cast_pe                 (cast_data_i_2_20),
    .ready_o_cast_pe                (cast_ready_o_2_20),
    .valid_o_cast_pe                (cast_valid_o_2_20),
    .data_o_cast_pe                 (cast_data_o_2_20),
    .ready_i_cast_pe                (cast_ready_i_2_20),

    .valid_i_merge_pe               (merge_valid_i_2_20),
    .data_i_merge_pe                (merge_data_i_2_20),
    .ready_o_merge_pe               (merge_ready_o_2_20),
    .valid_o_merge_pe               (merge_valid_o_2_20),
    .data_o_merge_pe                (merge_data_o_2_20),
    .ready_i_merge_pe               (merge_ready_i_2_20),

    .valid_i_gather_pe              (gather_valid_i_2_20),
    .data_i_gather_pe               (gather_data_i_2_20),
    .ready_o_gather_pe              (gather_ready_o_2_20),
    .valid_o_gather_pe              (gather_valid_o_2_20),
    .data_o_gather_pe               (gather_data_o_2_20),
    .ready_i_gather_pe              (gather_ready_i_2_20),

    .credit_upd                     (credit_upd[2][20])
);


network_interface #(
    .cast_out                       (cast_out_2_21),
    .gather_out                     (gather_out_2_21),
    .cast_sid                       (cast_sid_2_21),
    .gather_sid                     (gather_sid_2_21)
)ni_2_21(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[2][21]),
    .data_i_cast_nw                 (data_o_cast_nw[2][21]),
    .ready_o_cast_nw                (ready_i_cast_nw[2][21]),
    .valid_o_cast_nw                (valid_i_cast_nw[2][21]),
    .data_o_cast_nw                 (data_i_cast_nw[2][21]),
    .ready_i_cast_nw                (ready_o_cast_nw[2][21]),

    .valid_i_gather_nw              (valid_o_gather_nw[2][21]),
    .data_i_gather_nw               (data_o_gather_nw[2][21]),
    .ready_o_gather_nw              (ready_i_gather_nw[2][21]),
    .valid_o_gather_nw              (valid_i_gather_nw[2][21]),
    .data_o_gather_nw               (data_i_gather_nw[2][21]),
    .ready_i_gather_nw              (ready_o_gather_nw[2][21]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[2][21]),
    .data_i_merge_nw                (data_o_merge_nw[2][21]),
    .ready_o_merge_nw               (ready_i_merge_nw[2][21]),
    .valid_o_merge_nw               (valid_i_merge_nw[2][21]),
    .data_o_merge_nw                (data_i_merge_nw[2][21]),
    .ready_i_merge_nw               (ready_o_merge_nw[2][21]),

    .valid_i_cast_pe                (cast_valid_i_2_21),
    .data_i_cast_pe                 (cast_data_i_2_21),
    .ready_o_cast_pe                (cast_ready_o_2_21),
    .valid_o_cast_pe                (cast_valid_o_2_21),
    .data_o_cast_pe                 (cast_data_o_2_21),
    .ready_i_cast_pe                (cast_ready_i_2_21),

    .valid_i_merge_pe               (merge_valid_i_2_21),
    .data_i_merge_pe                (merge_data_i_2_21),
    .ready_o_merge_pe               (merge_ready_o_2_21),
    .valid_o_merge_pe               (merge_valid_o_2_21),
    .data_o_merge_pe                (merge_data_o_2_21),
    .ready_i_merge_pe               (merge_ready_i_2_21),

    .valid_i_gather_pe              (gather_valid_i_2_21),
    .data_i_gather_pe               (gather_data_i_2_21),
    .ready_o_gather_pe              (gather_ready_o_2_21),
    .valid_o_gather_pe              (gather_valid_o_2_21),
    .data_o_gather_pe               (gather_data_o_2_21),
    .ready_i_gather_pe              (gather_ready_i_2_21),

    .credit_upd                     (credit_upd[2][21])
);


network_interface #(
    .cast_out                       (cast_out_2_22),
    .gather_out                     (gather_out_2_22),
    .cast_sid                       (cast_sid_2_22),
    .gather_sid                     (gather_sid_2_22)
)ni_2_22(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[2][22]),
    .data_i_cast_nw                 (data_o_cast_nw[2][22]),
    .ready_o_cast_nw                (ready_i_cast_nw[2][22]),
    .valid_o_cast_nw                (valid_i_cast_nw[2][22]),
    .data_o_cast_nw                 (data_i_cast_nw[2][22]),
    .ready_i_cast_nw                (ready_o_cast_nw[2][22]),

    .valid_i_gather_nw              (valid_o_gather_nw[2][22]),
    .data_i_gather_nw               (data_o_gather_nw[2][22]),
    .ready_o_gather_nw              (ready_i_gather_nw[2][22]),
    .valid_o_gather_nw              (valid_i_gather_nw[2][22]),
    .data_o_gather_nw               (data_i_gather_nw[2][22]),
    .ready_i_gather_nw              (ready_o_gather_nw[2][22]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[2][22]),
    .data_i_merge_nw                (data_o_merge_nw[2][22]),
    .ready_o_merge_nw               (ready_i_merge_nw[2][22]),
    .valid_o_merge_nw               (valid_i_merge_nw[2][22]),
    .data_o_merge_nw                (data_i_merge_nw[2][22]),
    .ready_i_merge_nw               (ready_o_merge_nw[2][22]),

    .valid_i_cast_pe                (cast_valid_i_2_22),
    .data_i_cast_pe                 (cast_data_i_2_22),
    .ready_o_cast_pe                (cast_ready_o_2_22),
    .valid_o_cast_pe                (cast_valid_o_2_22),
    .data_o_cast_pe                 (cast_data_o_2_22),
    .ready_i_cast_pe                (cast_ready_i_2_22),

    .valid_i_merge_pe               (merge_valid_i_2_22),
    .data_i_merge_pe                (merge_data_i_2_22),
    .ready_o_merge_pe               (merge_ready_o_2_22),
    .valid_o_merge_pe               (merge_valid_o_2_22),
    .data_o_merge_pe                (merge_data_o_2_22),
    .ready_i_merge_pe               (merge_ready_i_2_22),

    .valid_i_gather_pe              (gather_valid_i_2_22),
    .data_i_gather_pe               (gather_data_i_2_22),
    .ready_o_gather_pe              (gather_ready_o_2_22),
    .valid_o_gather_pe              (gather_valid_o_2_22),
    .data_o_gather_pe               (gather_data_o_2_22),
    .ready_i_gather_pe              (gather_ready_i_2_22),

    .credit_upd                     (credit_upd[2][22])
);


network_interface #(
    .cast_out                       (cast_out_2_23),
    .gather_out                     (gather_out_2_23),
    .cast_sid                       (cast_sid_2_23),
    .gather_sid                     (gather_sid_2_23)
)ni_2_23(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[2][23]),
    .data_i_cast_nw                 (data_o_cast_nw[2][23]),
    .ready_o_cast_nw                (ready_i_cast_nw[2][23]),
    .valid_o_cast_nw                (valid_i_cast_nw[2][23]),
    .data_o_cast_nw                 (data_i_cast_nw[2][23]),
    .ready_i_cast_nw                (ready_o_cast_nw[2][23]),

    .valid_i_gather_nw              (valid_o_gather_nw[2][23]),
    .data_i_gather_nw               (data_o_gather_nw[2][23]),
    .ready_o_gather_nw              (ready_i_gather_nw[2][23]),
    .valid_o_gather_nw              (valid_i_gather_nw[2][23]),
    .data_o_gather_nw               (data_i_gather_nw[2][23]),
    .ready_i_gather_nw              (ready_o_gather_nw[2][23]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[2][23]),
    .data_i_merge_nw                (data_o_merge_nw[2][23]),
    .ready_o_merge_nw               (ready_i_merge_nw[2][23]),
    .valid_o_merge_nw               (valid_i_merge_nw[2][23]),
    .data_o_merge_nw                (data_i_merge_nw[2][23]),
    .ready_i_merge_nw               (ready_o_merge_nw[2][23]),

    .valid_i_cast_pe                (cast_valid_i_2_23),
    .data_i_cast_pe                 (cast_data_i_2_23),
    .ready_o_cast_pe                (cast_ready_o_2_23),
    .valid_o_cast_pe                (cast_valid_o_2_23),
    .data_o_cast_pe                 (cast_data_o_2_23),
    .ready_i_cast_pe                (cast_ready_i_2_23),

    .valid_i_merge_pe               (merge_valid_i_2_23),
    .data_i_merge_pe                (merge_data_i_2_23),
    .ready_o_merge_pe               (merge_ready_o_2_23),
    .valid_o_merge_pe               (merge_valid_o_2_23),
    .data_o_merge_pe                (merge_data_o_2_23),
    .ready_i_merge_pe               (merge_ready_i_2_23),

    .valid_i_gather_pe              (gather_valid_i_2_23),
    .data_i_gather_pe               (gather_data_i_2_23),
    .ready_o_gather_pe              (gather_ready_o_2_23),
    .valid_o_gather_pe              (gather_valid_o_2_23),
    .data_o_gather_pe               (gather_data_o_2_23),
    .ready_i_gather_pe              (gather_ready_i_2_23),

    .credit_upd                     (credit_upd[2][23])
);


network_interface #(
    .cast_out                       (cast_out_2_24),
    .gather_out                     (gather_out_2_24),
    .cast_sid                       (cast_sid_2_24),
    .gather_sid                     (gather_sid_2_24)
)ni_2_24(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[2][24]),
    .data_i_cast_nw                 (data_o_cast_nw[2][24]),
    .ready_o_cast_nw                (ready_i_cast_nw[2][24]),
    .valid_o_cast_nw                (valid_i_cast_nw[2][24]),
    .data_o_cast_nw                 (data_i_cast_nw[2][24]),
    .ready_i_cast_nw                (ready_o_cast_nw[2][24]),

    .valid_i_gather_nw              (valid_o_gather_nw[2][24]),
    .data_i_gather_nw               (data_o_gather_nw[2][24]),
    .ready_o_gather_nw              (ready_i_gather_nw[2][24]),
    .valid_o_gather_nw              (valid_i_gather_nw[2][24]),
    .data_o_gather_nw               (data_i_gather_nw[2][24]),
    .ready_i_gather_nw              (ready_o_gather_nw[2][24]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[2][24]),
    .data_i_merge_nw                (data_o_merge_nw[2][24]),
    .ready_o_merge_nw               (ready_i_merge_nw[2][24]),
    .valid_o_merge_nw               (valid_i_merge_nw[2][24]),
    .data_o_merge_nw                (data_i_merge_nw[2][24]),
    .ready_i_merge_nw               (ready_o_merge_nw[2][24]),

    .valid_i_cast_pe                (cast_valid_i_2_24),
    .data_i_cast_pe                 (cast_data_i_2_24),
    .ready_o_cast_pe                (cast_ready_o_2_24),
    .valid_o_cast_pe                (cast_valid_o_2_24),
    .data_o_cast_pe                 (cast_data_o_2_24),
    .ready_i_cast_pe                (cast_ready_i_2_24),

    .valid_i_merge_pe               (merge_valid_i_2_24),
    .data_i_merge_pe                (merge_data_i_2_24),
    .ready_o_merge_pe               (merge_ready_o_2_24),
    .valid_o_merge_pe               (merge_valid_o_2_24),
    .data_o_merge_pe                (merge_data_o_2_24),
    .ready_i_merge_pe               (merge_ready_i_2_24),

    .valid_i_gather_pe              (gather_valid_i_2_24),
    .data_i_gather_pe               (gather_data_i_2_24),
    .ready_o_gather_pe              (gather_ready_o_2_24),
    .valid_o_gather_pe              (gather_valid_o_2_24),
    .data_o_gather_pe               (gather_data_o_2_24),
    .ready_i_gather_pe              (gather_ready_i_2_24),

    .credit_upd                     (credit_upd[2][24])
);


network_interface #(
    .cast_out                       (cast_out_3_0),
    .gather_out                     (gather_out_3_0),
    .cast_sid                       (cast_sid_3_0),
    .gather_sid                     (gather_sid_3_0)
)ni_3_0(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[3][0]),
    .data_i_cast_nw                 (data_o_cast_nw[3][0]),
    .ready_o_cast_nw                (ready_i_cast_nw[3][0]),
    .valid_o_cast_nw                (valid_i_cast_nw[3][0]),
    .data_o_cast_nw                 (data_i_cast_nw[3][0]),
    .ready_i_cast_nw                (ready_o_cast_nw[3][0]),

    .valid_i_gather_nw              (valid_o_gather_nw[3][0]),
    .data_i_gather_nw               (data_o_gather_nw[3][0]),
    .ready_o_gather_nw              (ready_i_gather_nw[3][0]),
    .valid_o_gather_nw              (valid_i_gather_nw[3][0]),
    .data_o_gather_nw               (data_i_gather_nw[3][0]),
    .ready_i_gather_nw              (ready_o_gather_nw[3][0]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[3][0]),
    .data_i_merge_nw                (data_o_merge_nw[3][0]),
    .ready_o_merge_nw               (ready_i_merge_nw[3][0]),
    .valid_o_merge_nw               (valid_i_merge_nw[3][0]),
    .data_o_merge_nw                (data_i_merge_nw[3][0]),
    .ready_i_merge_nw               (ready_o_merge_nw[3][0]),

    .valid_i_cast_pe                (cast_valid_i_3_0),
    .data_i_cast_pe                 (cast_data_i_3_0),
    .ready_o_cast_pe                (cast_ready_o_3_0),
    .valid_o_cast_pe                (cast_valid_o_3_0),
    .data_o_cast_pe                 (cast_data_o_3_0),
    .ready_i_cast_pe                (cast_ready_i_3_0),

    .valid_i_merge_pe               (merge_valid_i_3_0),
    .data_i_merge_pe                (merge_data_i_3_0),
    .ready_o_merge_pe               (merge_ready_o_3_0),
    .valid_o_merge_pe               (merge_valid_o_3_0),
    .data_o_merge_pe                (merge_data_o_3_0),
    .ready_i_merge_pe               (merge_ready_i_3_0),

    .valid_i_gather_pe              (gather_valid_i_3_0),
    .data_i_gather_pe               (gather_data_i_3_0),
    .ready_o_gather_pe              (gather_ready_o_3_0),
    .valid_o_gather_pe              (gather_valid_o_3_0),
    .data_o_gather_pe               (gather_data_o_3_0),
    .ready_i_gather_pe              (gather_ready_i_3_0),

    .credit_upd                     (credit_upd[3][0])
);


network_interface #(
    .cast_out                       (cast_out_3_1),
    .gather_out                     (gather_out_3_1),
    .cast_sid                       (cast_sid_3_1),
    .gather_sid                     (gather_sid_3_1)
)ni_3_1(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[3][1]),
    .data_i_cast_nw                 (data_o_cast_nw[3][1]),
    .ready_o_cast_nw                (ready_i_cast_nw[3][1]),
    .valid_o_cast_nw                (valid_i_cast_nw[3][1]),
    .data_o_cast_nw                 (data_i_cast_nw[3][1]),
    .ready_i_cast_nw                (ready_o_cast_nw[3][1]),

    .valid_i_gather_nw              (valid_o_gather_nw[3][1]),
    .data_i_gather_nw               (data_o_gather_nw[3][1]),
    .ready_o_gather_nw              (ready_i_gather_nw[3][1]),
    .valid_o_gather_nw              (valid_i_gather_nw[3][1]),
    .data_o_gather_nw               (data_i_gather_nw[3][1]),
    .ready_i_gather_nw              (ready_o_gather_nw[3][1]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[3][1]),
    .data_i_merge_nw                (data_o_merge_nw[3][1]),
    .ready_o_merge_nw               (ready_i_merge_nw[3][1]),
    .valid_o_merge_nw               (valid_i_merge_nw[3][1]),
    .data_o_merge_nw                (data_i_merge_nw[3][1]),
    .ready_i_merge_nw               (ready_o_merge_nw[3][1]),

    .valid_i_cast_pe                (cast_valid_i_3_1),
    .data_i_cast_pe                 (cast_data_i_3_1),
    .ready_o_cast_pe                (cast_ready_o_3_1),
    .valid_o_cast_pe                (cast_valid_o_3_1),
    .data_o_cast_pe                 (cast_data_o_3_1),
    .ready_i_cast_pe                (cast_ready_i_3_1),

    .valid_i_merge_pe               (merge_valid_i_3_1),
    .data_i_merge_pe                (merge_data_i_3_1),
    .ready_o_merge_pe               (merge_ready_o_3_1),
    .valid_o_merge_pe               (merge_valid_o_3_1),
    .data_o_merge_pe                (merge_data_o_3_1),
    .ready_i_merge_pe               (merge_ready_i_3_1),

    .valid_i_gather_pe              (gather_valid_i_3_1),
    .data_i_gather_pe               (gather_data_i_3_1),
    .ready_o_gather_pe              (gather_ready_o_3_1),
    .valid_o_gather_pe              (gather_valid_o_3_1),
    .data_o_gather_pe               (gather_data_o_3_1),
    .ready_i_gather_pe              (gather_ready_i_3_1),

    .credit_upd                     (credit_upd[3][1])
);


network_interface #(
    .cast_out                       (cast_out_3_2),
    .gather_out                     (gather_out_3_2),
    .cast_sid                       (cast_sid_3_2),
    .gather_sid                     (gather_sid_3_2)
)ni_3_2(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[3][2]),
    .data_i_cast_nw                 (data_o_cast_nw[3][2]),
    .ready_o_cast_nw                (ready_i_cast_nw[3][2]),
    .valid_o_cast_nw                (valid_i_cast_nw[3][2]),
    .data_o_cast_nw                 (data_i_cast_nw[3][2]),
    .ready_i_cast_nw                (ready_o_cast_nw[3][2]),

    .valid_i_gather_nw              (valid_o_gather_nw[3][2]),
    .data_i_gather_nw               (data_o_gather_nw[3][2]),
    .ready_o_gather_nw              (ready_i_gather_nw[3][2]),
    .valid_o_gather_nw              (valid_i_gather_nw[3][2]),
    .data_o_gather_nw               (data_i_gather_nw[3][2]),
    .ready_i_gather_nw              (ready_o_gather_nw[3][2]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[3][2]),
    .data_i_merge_nw                (data_o_merge_nw[3][2]),
    .ready_o_merge_nw               (ready_i_merge_nw[3][2]),
    .valid_o_merge_nw               (valid_i_merge_nw[3][2]),
    .data_o_merge_nw                (data_i_merge_nw[3][2]),
    .ready_i_merge_nw               (ready_o_merge_nw[3][2]),

    .valid_i_cast_pe                (cast_valid_i_3_2),
    .data_i_cast_pe                 (cast_data_i_3_2),
    .ready_o_cast_pe                (cast_ready_o_3_2),
    .valid_o_cast_pe                (cast_valid_o_3_2),
    .data_o_cast_pe                 (cast_data_o_3_2),
    .ready_i_cast_pe                (cast_ready_i_3_2),

    .valid_i_merge_pe               (merge_valid_i_3_2),
    .data_i_merge_pe                (merge_data_i_3_2),
    .ready_o_merge_pe               (merge_ready_o_3_2),
    .valid_o_merge_pe               (merge_valid_o_3_2),
    .data_o_merge_pe                (merge_data_o_3_2),
    .ready_i_merge_pe               (merge_ready_i_3_2),

    .valid_i_gather_pe              (gather_valid_i_3_2),
    .data_i_gather_pe               (gather_data_i_3_2),
    .ready_o_gather_pe              (gather_ready_o_3_2),
    .valid_o_gather_pe              (gather_valid_o_3_2),
    .data_o_gather_pe               (gather_data_o_3_2),
    .ready_i_gather_pe              (gather_ready_i_3_2),

    .credit_upd                     (credit_upd[3][2])
);


network_interface #(
    .cast_out                       (cast_out_3_3),
    .gather_out                     (gather_out_3_3),
    .cast_sid                       (cast_sid_3_3),
    .gather_sid                     (gather_sid_3_3)
)ni_3_3(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[3][3]),
    .data_i_cast_nw                 (data_o_cast_nw[3][3]),
    .ready_o_cast_nw                (ready_i_cast_nw[3][3]),
    .valid_o_cast_nw                (valid_i_cast_nw[3][3]),
    .data_o_cast_nw                 (data_i_cast_nw[3][3]),
    .ready_i_cast_nw                (ready_o_cast_nw[3][3]),

    .valid_i_gather_nw              (valid_o_gather_nw[3][3]),
    .data_i_gather_nw               (data_o_gather_nw[3][3]),
    .ready_o_gather_nw              (ready_i_gather_nw[3][3]),
    .valid_o_gather_nw              (valid_i_gather_nw[3][3]),
    .data_o_gather_nw               (data_i_gather_nw[3][3]),
    .ready_i_gather_nw              (ready_o_gather_nw[3][3]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[3][3]),
    .data_i_merge_nw                (data_o_merge_nw[3][3]),
    .ready_o_merge_nw               (ready_i_merge_nw[3][3]),
    .valid_o_merge_nw               (valid_i_merge_nw[3][3]),
    .data_o_merge_nw                (data_i_merge_nw[3][3]),
    .ready_i_merge_nw               (ready_o_merge_nw[3][3]),

    .valid_i_cast_pe                (cast_valid_i_3_3),
    .data_i_cast_pe                 (cast_data_i_3_3),
    .ready_o_cast_pe                (cast_ready_o_3_3),
    .valid_o_cast_pe                (cast_valid_o_3_3),
    .data_o_cast_pe                 (cast_data_o_3_3),
    .ready_i_cast_pe                (cast_ready_i_3_3),

    .valid_i_merge_pe               (merge_valid_i_3_3),
    .data_i_merge_pe                (merge_data_i_3_3),
    .ready_o_merge_pe               (merge_ready_o_3_3),
    .valid_o_merge_pe               (merge_valid_o_3_3),
    .data_o_merge_pe                (merge_data_o_3_3),
    .ready_i_merge_pe               (merge_ready_i_3_3),

    .valid_i_gather_pe              (gather_valid_i_3_3),
    .data_i_gather_pe               (gather_data_i_3_3),
    .ready_o_gather_pe              (gather_ready_o_3_3),
    .valid_o_gather_pe              (gather_valid_o_3_3),
    .data_o_gather_pe               (gather_data_o_3_3),
    .ready_i_gather_pe              (gather_ready_i_3_3),

    .credit_upd                     (credit_upd[3][3])
);


network_interface #(
    .cast_out                       (cast_out_3_4),
    .gather_out                     (gather_out_3_4),
    .cast_sid                       (cast_sid_3_4),
    .gather_sid                     (gather_sid_3_4)
)ni_3_4(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[3][4]),
    .data_i_cast_nw                 (data_o_cast_nw[3][4]),
    .ready_o_cast_nw                (ready_i_cast_nw[3][4]),
    .valid_o_cast_nw                (valid_i_cast_nw[3][4]),
    .data_o_cast_nw                 (data_i_cast_nw[3][4]),
    .ready_i_cast_nw                (ready_o_cast_nw[3][4]),

    .valid_i_gather_nw              (valid_o_gather_nw[3][4]),
    .data_i_gather_nw               (data_o_gather_nw[3][4]),
    .ready_o_gather_nw              (ready_i_gather_nw[3][4]),
    .valid_o_gather_nw              (valid_i_gather_nw[3][4]),
    .data_o_gather_nw               (data_i_gather_nw[3][4]),
    .ready_i_gather_nw              (ready_o_gather_nw[3][4]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[3][4]),
    .data_i_merge_nw                (data_o_merge_nw[3][4]),
    .ready_o_merge_nw               (ready_i_merge_nw[3][4]),
    .valid_o_merge_nw               (valid_i_merge_nw[3][4]),
    .data_o_merge_nw                (data_i_merge_nw[3][4]),
    .ready_i_merge_nw               (ready_o_merge_nw[3][4]),

    .valid_i_cast_pe                (cast_valid_i_3_4),
    .data_i_cast_pe                 (cast_data_i_3_4),
    .ready_o_cast_pe                (cast_ready_o_3_4),
    .valid_o_cast_pe                (cast_valid_o_3_4),
    .data_o_cast_pe                 (cast_data_o_3_4),
    .ready_i_cast_pe                (cast_ready_i_3_4),

    .valid_i_merge_pe               (merge_valid_i_3_4),
    .data_i_merge_pe                (merge_data_i_3_4),
    .ready_o_merge_pe               (merge_ready_o_3_4),
    .valid_o_merge_pe               (merge_valid_o_3_4),
    .data_o_merge_pe                (merge_data_o_3_4),
    .ready_i_merge_pe               (merge_ready_i_3_4),

    .valid_i_gather_pe              (gather_valid_i_3_4),
    .data_i_gather_pe               (gather_data_i_3_4),
    .ready_o_gather_pe              (gather_ready_o_3_4),
    .valid_o_gather_pe              (gather_valid_o_3_4),
    .data_o_gather_pe               (gather_data_o_3_4),
    .ready_i_gather_pe              (gather_ready_i_3_4),

    .credit_upd                     (credit_upd[3][4])
);


network_interface #(
    .cast_out                       (cast_out_3_5),
    .gather_out                     (gather_out_3_5),
    .cast_sid                       (cast_sid_3_5),
    .gather_sid                     (gather_sid_3_5)
)ni_3_5(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[3][5]),
    .data_i_cast_nw                 (data_o_cast_nw[3][5]),
    .ready_o_cast_nw                (ready_i_cast_nw[3][5]),
    .valid_o_cast_nw                (valid_i_cast_nw[3][5]),
    .data_o_cast_nw                 (data_i_cast_nw[3][5]),
    .ready_i_cast_nw                (ready_o_cast_nw[3][5]),

    .valid_i_gather_nw              (valid_o_gather_nw[3][5]),
    .data_i_gather_nw               (data_o_gather_nw[3][5]),
    .ready_o_gather_nw              (ready_i_gather_nw[3][5]),
    .valid_o_gather_nw              (valid_i_gather_nw[3][5]),
    .data_o_gather_nw               (data_i_gather_nw[3][5]),
    .ready_i_gather_nw              (ready_o_gather_nw[3][5]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[3][5]),
    .data_i_merge_nw                (data_o_merge_nw[3][5]),
    .ready_o_merge_nw               (ready_i_merge_nw[3][5]),
    .valid_o_merge_nw               (valid_i_merge_nw[3][5]),
    .data_o_merge_nw                (data_i_merge_nw[3][5]),
    .ready_i_merge_nw               (ready_o_merge_nw[3][5]),

    .valid_i_cast_pe                (cast_valid_i_3_5),
    .data_i_cast_pe                 (cast_data_i_3_5),
    .ready_o_cast_pe                (cast_ready_o_3_5),
    .valid_o_cast_pe                (cast_valid_o_3_5),
    .data_o_cast_pe                 (cast_data_o_3_5),
    .ready_i_cast_pe                (cast_ready_i_3_5),

    .valid_i_merge_pe               (merge_valid_i_3_5),
    .data_i_merge_pe                (merge_data_i_3_5),
    .ready_o_merge_pe               (merge_ready_o_3_5),
    .valid_o_merge_pe               (merge_valid_o_3_5),
    .data_o_merge_pe                (merge_data_o_3_5),
    .ready_i_merge_pe               (merge_ready_i_3_5),

    .valid_i_gather_pe              (gather_valid_i_3_5),
    .data_i_gather_pe               (gather_data_i_3_5),
    .ready_o_gather_pe              (gather_ready_o_3_5),
    .valid_o_gather_pe              (gather_valid_o_3_5),
    .data_o_gather_pe               (gather_data_o_3_5),
    .ready_i_gather_pe              (gather_ready_i_3_5),

    .credit_upd                     (credit_upd[3][5])
);


network_interface #(
    .cast_out                       (cast_out_3_6),
    .gather_out                     (gather_out_3_6),
    .cast_sid                       (cast_sid_3_6),
    .gather_sid                     (gather_sid_3_6)
)ni_3_6(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[3][6]),
    .data_i_cast_nw                 (data_o_cast_nw[3][6]),
    .ready_o_cast_nw                (ready_i_cast_nw[3][6]),
    .valid_o_cast_nw                (valid_i_cast_nw[3][6]),
    .data_o_cast_nw                 (data_i_cast_nw[3][6]),
    .ready_i_cast_nw                (ready_o_cast_nw[3][6]),

    .valid_i_gather_nw              (valid_o_gather_nw[3][6]),
    .data_i_gather_nw               (data_o_gather_nw[3][6]),
    .ready_o_gather_nw              (ready_i_gather_nw[3][6]),
    .valid_o_gather_nw              (valid_i_gather_nw[3][6]),
    .data_o_gather_nw               (data_i_gather_nw[3][6]),
    .ready_i_gather_nw              (ready_o_gather_nw[3][6]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[3][6]),
    .data_i_merge_nw                (data_o_merge_nw[3][6]),
    .ready_o_merge_nw               (ready_i_merge_nw[3][6]),
    .valid_o_merge_nw               (valid_i_merge_nw[3][6]),
    .data_o_merge_nw                (data_i_merge_nw[3][6]),
    .ready_i_merge_nw               (ready_o_merge_nw[3][6]),

    .valid_i_cast_pe                (cast_valid_i_3_6),
    .data_i_cast_pe                 (cast_data_i_3_6),
    .ready_o_cast_pe                (cast_ready_o_3_6),
    .valid_o_cast_pe                (cast_valid_o_3_6),
    .data_o_cast_pe                 (cast_data_o_3_6),
    .ready_i_cast_pe                (cast_ready_i_3_6),

    .valid_i_merge_pe               (merge_valid_i_3_6),
    .data_i_merge_pe                (merge_data_i_3_6),
    .ready_o_merge_pe               (merge_ready_o_3_6),
    .valid_o_merge_pe               (merge_valid_o_3_6),
    .data_o_merge_pe                (merge_data_o_3_6),
    .ready_i_merge_pe               (merge_ready_i_3_6),

    .valid_i_gather_pe              (gather_valid_i_3_6),
    .data_i_gather_pe               (gather_data_i_3_6),
    .ready_o_gather_pe              (gather_ready_o_3_6),
    .valid_o_gather_pe              (gather_valid_o_3_6),
    .data_o_gather_pe               (gather_data_o_3_6),
    .ready_i_gather_pe              (gather_ready_i_3_6),

    .credit_upd                     (credit_upd[3][6])
);


network_interface #(
    .cast_out                       (cast_out_3_7),
    .gather_out                     (gather_out_3_7),
    .cast_sid                       (cast_sid_3_7),
    .gather_sid                     (gather_sid_3_7)
)ni_3_7(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[3][7]),
    .data_i_cast_nw                 (data_o_cast_nw[3][7]),
    .ready_o_cast_nw                (ready_i_cast_nw[3][7]),
    .valid_o_cast_nw                (valid_i_cast_nw[3][7]),
    .data_o_cast_nw                 (data_i_cast_nw[3][7]),
    .ready_i_cast_nw                (ready_o_cast_nw[3][7]),

    .valid_i_gather_nw              (valid_o_gather_nw[3][7]),
    .data_i_gather_nw               (data_o_gather_nw[3][7]),
    .ready_o_gather_nw              (ready_i_gather_nw[3][7]),
    .valid_o_gather_nw              (valid_i_gather_nw[3][7]),
    .data_o_gather_nw               (data_i_gather_nw[3][7]),
    .ready_i_gather_nw              (ready_o_gather_nw[3][7]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[3][7]),
    .data_i_merge_nw                (data_o_merge_nw[3][7]),
    .ready_o_merge_nw               (ready_i_merge_nw[3][7]),
    .valid_o_merge_nw               (valid_i_merge_nw[3][7]),
    .data_o_merge_nw                (data_i_merge_nw[3][7]),
    .ready_i_merge_nw               (ready_o_merge_nw[3][7]),

    .valid_i_cast_pe                (cast_valid_i_3_7),
    .data_i_cast_pe                 (cast_data_i_3_7),
    .ready_o_cast_pe                (cast_ready_o_3_7),
    .valid_o_cast_pe                (cast_valid_o_3_7),
    .data_o_cast_pe                 (cast_data_o_3_7),
    .ready_i_cast_pe                (cast_ready_i_3_7),

    .valid_i_merge_pe               (merge_valid_i_3_7),
    .data_i_merge_pe                (merge_data_i_3_7),
    .ready_o_merge_pe               (merge_ready_o_3_7),
    .valid_o_merge_pe               (merge_valid_o_3_7),
    .data_o_merge_pe                (merge_data_o_3_7),
    .ready_i_merge_pe               (merge_ready_i_3_7),

    .valid_i_gather_pe              (gather_valid_i_3_7),
    .data_i_gather_pe               (gather_data_i_3_7),
    .ready_o_gather_pe              (gather_ready_o_3_7),
    .valid_o_gather_pe              (gather_valid_o_3_7),
    .data_o_gather_pe               (gather_data_o_3_7),
    .ready_i_gather_pe              (gather_ready_i_3_7),

    .credit_upd                     (credit_upd[3][7])
);


network_interface #(
    .cast_out                       (cast_out_3_8),
    .gather_out                     (gather_out_3_8),
    .cast_sid                       (cast_sid_3_8),
    .gather_sid                     (gather_sid_3_8)
)ni_3_8(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[3][8]),
    .data_i_cast_nw                 (data_o_cast_nw[3][8]),
    .ready_o_cast_nw                (ready_i_cast_nw[3][8]),
    .valid_o_cast_nw                (valid_i_cast_nw[3][8]),
    .data_o_cast_nw                 (data_i_cast_nw[3][8]),
    .ready_i_cast_nw                (ready_o_cast_nw[3][8]),

    .valid_i_gather_nw              (valid_o_gather_nw[3][8]),
    .data_i_gather_nw               (data_o_gather_nw[3][8]),
    .ready_o_gather_nw              (ready_i_gather_nw[3][8]),
    .valid_o_gather_nw              (valid_i_gather_nw[3][8]),
    .data_o_gather_nw               (data_i_gather_nw[3][8]),
    .ready_i_gather_nw              (ready_o_gather_nw[3][8]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[3][8]),
    .data_i_merge_nw                (data_o_merge_nw[3][8]),
    .ready_o_merge_nw               (ready_i_merge_nw[3][8]),
    .valid_o_merge_nw               (valid_i_merge_nw[3][8]),
    .data_o_merge_nw                (data_i_merge_nw[3][8]),
    .ready_i_merge_nw               (ready_o_merge_nw[3][8]),

    .valid_i_cast_pe                (cast_valid_i_3_8),
    .data_i_cast_pe                 (cast_data_i_3_8),
    .ready_o_cast_pe                (cast_ready_o_3_8),
    .valid_o_cast_pe                (cast_valid_o_3_8),
    .data_o_cast_pe                 (cast_data_o_3_8),
    .ready_i_cast_pe                (cast_ready_i_3_8),

    .valid_i_merge_pe               (merge_valid_i_3_8),
    .data_i_merge_pe                (merge_data_i_3_8),
    .ready_o_merge_pe               (merge_ready_o_3_8),
    .valid_o_merge_pe               (merge_valid_o_3_8),
    .data_o_merge_pe                (merge_data_o_3_8),
    .ready_i_merge_pe               (merge_ready_i_3_8),

    .valid_i_gather_pe              (gather_valid_i_3_8),
    .data_i_gather_pe               (gather_data_i_3_8),
    .ready_o_gather_pe              (gather_ready_o_3_8),
    .valid_o_gather_pe              (gather_valid_o_3_8),
    .data_o_gather_pe               (gather_data_o_3_8),
    .ready_i_gather_pe              (gather_ready_i_3_8),

    .credit_upd                     (credit_upd[3][8])
);


network_interface #(
    .cast_out                       (cast_out_3_9),
    .gather_out                     (gather_out_3_9),
    .cast_sid                       (cast_sid_3_9),
    .gather_sid                     (gather_sid_3_9)
)ni_3_9(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[3][9]),
    .data_i_cast_nw                 (data_o_cast_nw[3][9]),
    .ready_o_cast_nw                (ready_i_cast_nw[3][9]),
    .valid_o_cast_nw                (valid_i_cast_nw[3][9]),
    .data_o_cast_nw                 (data_i_cast_nw[3][9]),
    .ready_i_cast_nw                (ready_o_cast_nw[3][9]),

    .valid_i_gather_nw              (valid_o_gather_nw[3][9]),
    .data_i_gather_nw               (data_o_gather_nw[3][9]),
    .ready_o_gather_nw              (ready_i_gather_nw[3][9]),
    .valid_o_gather_nw              (valid_i_gather_nw[3][9]),
    .data_o_gather_nw               (data_i_gather_nw[3][9]),
    .ready_i_gather_nw              (ready_o_gather_nw[3][9]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[3][9]),
    .data_i_merge_nw                (data_o_merge_nw[3][9]),
    .ready_o_merge_nw               (ready_i_merge_nw[3][9]),
    .valid_o_merge_nw               (valid_i_merge_nw[3][9]),
    .data_o_merge_nw                (data_i_merge_nw[3][9]),
    .ready_i_merge_nw               (ready_o_merge_nw[3][9]),

    .valid_i_cast_pe                (cast_valid_i_3_9),
    .data_i_cast_pe                 (cast_data_i_3_9),
    .ready_o_cast_pe                (cast_ready_o_3_9),
    .valid_o_cast_pe                (cast_valid_o_3_9),
    .data_o_cast_pe                 (cast_data_o_3_9),
    .ready_i_cast_pe                (cast_ready_i_3_9),

    .valid_i_merge_pe               (merge_valid_i_3_9),
    .data_i_merge_pe                (merge_data_i_3_9),
    .ready_o_merge_pe               (merge_ready_o_3_9),
    .valid_o_merge_pe               (merge_valid_o_3_9),
    .data_o_merge_pe                (merge_data_o_3_9),
    .ready_i_merge_pe               (merge_ready_i_3_9),

    .valid_i_gather_pe              (gather_valid_i_3_9),
    .data_i_gather_pe               (gather_data_i_3_9),
    .ready_o_gather_pe              (gather_ready_o_3_9),
    .valid_o_gather_pe              (gather_valid_o_3_9),
    .data_o_gather_pe               (gather_data_o_3_9),
    .ready_i_gather_pe              (gather_ready_i_3_9),

    .credit_upd                     (credit_upd[3][9])
);


network_interface #(
    .cast_out                       (cast_out_3_10),
    .gather_out                     (gather_out_3_10),
    .cast_sid                       (cast_sid_3_10),
    .gather_sid                     (gather_sid_3_10)
)ni_3_10(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[3][10]),
    .data_i_cast_nw                 (data_o_cast_nw[3][10]),
    .ready_o_cast_nw                (ready_i_cast_nw[3][10]),
    .valid_o_cast_nw                (valid_i_cast_nw[3][10]),
    .data_o_cast_nw                 (data_i_cast_nw[3][10]),
    .ready_i_cast_nw                (ready_o_cast_nw[3][10]),

    .valid_i_gather_nw              (valid_o_gather_nw[3][10]),
    .data_i_gather_nw               (data_o_gather_nw[3][10]),
    .ready_o_gather_nw              (ready_i_gather_nw[3][10]),
    .valid_o_gather_nw              (valid_i_gather_nw[3][10]),
    .data_o_gather_nw               (data_i_gather_nw[3][10]),
    .ready_i_gather_nw              (ready_o_gather_nw[3][10]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[3][10]),
    .data_i_merge_nw                (data_o_merge_nw[3][10]),
    .ready_o_merge_nw               (ready_i_merge_nw[3][10]),
    .valid_o_merge_nw               (valid_i_merge_nw[3][10]),
    .data_o_merge_nw                (data_i_merge_nw[3][10]),
    .ready_i_merge_nw               (ready_o_merge_nw[3][10]),

    .valid_i_cast_pe                (cast_valid_i_3_10),
    .data_i_cast_pe                 (cast_data_i_3_10),
    .ready_o_cast_pe                (cast_ready_o_3_10),
    .valid_o_cast_pe                (cast_valid_o_3_10),
    .data_o_cast_pe                 (cast_data_o_3_10),
    .ready_i_cast_pe                (cast_ready_i_3_10),

    .valid_i_merge_pe               (merge_valid_i_3_10),
    .data_i_merge_pe                (merge_data_i_3_10),
    .ready_o_merge_pe               (merge_ready_o_3_10),
    .valid_o_merge_pe               (merge_valid_o_3_10),
    .data_o_merge_pe                (merge_data_o_3_10),
    .ready_i_merge_pe               (merge_ready_i_3_10),

    .valid_i_gather_pe              (gather_valid_i_3_10),
    .data_i_gather_pe               (gather_data_i_3_10),
    .ready_o_gather_pe              (gather_ready_o_3_10),
    .valid_o_gather_pe              (gather_valid_o_3_10),
    .data_o_gather_pe               (gather_data_o_3_10),
    .ready_i_gather_pe              (gather_ready_i_3_10),

    .credit_upd                     (credit_upd[3][10])
);


network_interface #(
    .cast_out                       (cast_out_3_11),
    .gather_out                     (gather_out_3_11),
    .cast_sid                       (cast_sid_3_11),
    .gather_sid                     (gather_sid_3_11)
)ni_3_11(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[3][11]),
    .data_i_cast_nw                 (data_o_cast_nw[3][11]),
    .ready_o_cast_nw                (ready_i_cast_nw[3][11]),
    .valid_o_cast_nw                (valid_i_cast_nw[3][11]),
    .data_o_cast_nw                 (data_i_cast_nw[3][11]),
    .ready_i_cast_nw                (ready_o_cast_nw[3][11]),

    .valid_i_gather_nw              (valid_o_gather_nw[3][11]),
    .data_i_gather_nw               (data_o_gather_nw[3][11]),
    .ready_o_gather_nw              (ready_i_gather_nw[3][11]),
    .valid_o_gather_nw              (valid_i_gather_nw[3][11]),
    .data_o_gather_nw               (data_i_gather_nw[3][11]),
    .ready_i_gather_nw              (ready_o_gather_nw[3][11]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[3][11]),
    .data_i_merge_nw                (data_o_merge_nw[3][11]),
    .ready_o_merge_nw               (ready_i_merge_nw[3][11]),
    .valid_o_merge_nw               (valid_i_merge_nw[3][11]),
    .data_o_merge_nw                (data_i_merge_nw[3][11]),
    .ready_i_merge_nw               (ready_o_merge_nw[3][11]),

    .valid_i_cast_pe                (cast_valid_i_3_11),
    .data_i_cast_pe                 (cast_data_i_3_11),
    .ready_o_cast_pe                (cast_ready_o_3_11),
    .valid_o_cast_pe                (cast_valid_o_3_11),
    .data_o_cast_pe                 (cast_data_o_3_11),
    .ready_i_cast_pe                (cast_ready_i_3_11),

    .valid_i_merge_pe               (merge_valid_i_3_11),
    .data_i_merge_pe                (merge_data_i_3_11),
    .ready_o_merge_pe               (merge_ready_o_3_11),
    .valid_o_merge_pe               (merge_valid_o_3_11),
    .data_o_merge_pe                (merge_data_o_3_11),
    .ready_i_merge_pe               (merge_ready_i_3_11),

    .valid_i_gather_pe              (gather_valid_i_3_11),
    .data_i_gather_pe               (gather_data_i_3_11),
    .ready_o_gather_pe              (gather_ready_o_3_11),
    .valid_o_gather_pe              (gather_valid_o_3_11),
    .data_o_gather_pe               (gather_data_o_3_11),
    .ready_i_gather_pe              (gather_ready_i_3_11),

    .credit_upd                     (credit_upd[3][11])
);


network_interface #(
    .cast_out                       (cast_out_3_12),
    .gather_out                     (gather_out_3_12),
    .cast_sid                       (cast_sid_3_12),
    .gather_sid                     (gather_sid_3_12)
)ni_3_12(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[3][12]),
    .data_i_cast_nw                 (data_o_cast_nw[3][12]),
    .ready_o_cast_nw                (ready_i_cast_nw[3][12]),
    .valid_o_cast_nw                (valid_i_cast_nw[3][12]),
    .data_o_cast_nw                 (data_i_cast_nw[3][12]),
    .ready_i_cast_nw                (ready_o_cast_nw[3][12]),

    .valid_i_gather_nw              (valid_o_gather_nw[3][12]),
    .data_i_gather_nw               (data_o_gather_nw[3][12]),
    .ready_o_gather_nw              (ready_i_gather_nw[3][12]),
    .valid_o_gather_nw              (valid_i_gather_nw[3][12]),
    .data_o_gather_nw               (data_i_gather_nw[3][12]),
    .ready_i_gather_nw              (ready_o_gather_nw[3][12]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[3][12]),
    .data_i_merge_nw                (data_o_merge_nw[3][12]),
    .ready_o_merge_nw               (ready_i_merge_nw[3][12]),
    .valid_o_merge_nw               (valid_i_merge_nw[3][12]),
    .data_o_merge_nw                (data_i_merge_nw[3][12]),
    .ready_i_merge_nw               (ready_o_merge_nw[3][12]),

    .valid_i_cast_pe                (cast_valid_i_3_12),
    .data_i_cast_pe                 (cast_data_i_3_12),
    .ready_o_cast_pe                (cast_ready_o_3_12),
    .valid_o_cast_pe                (cast_valid_o_3_12),
    .data_o_cast_pe                 (cast_data_o_3_12),
    .ready_i_cast_pe                (cast_ready_i_3_12),

    .valid_i_merge_pe               (merge_valid_i_3_12),
    .data_i_merge_pe                (merge_data_i_3_12),
    .ready_o_merge_pe               (merge_ready_o_3_12),
    .valid_o_merge_pe               (merge_valid_o_3_12),
    .data_o_merge_pe                (merge_data_o_3_12),
    .ready_i_merge_pe               (merge_ready_i_3_12),

    .valid_i_gather_pe              (gather_valid_i_3_12),
    .data_i_gather_pe               (gather_data_i_3_12),
    .ready_o_gather_pe              (gather_ready_o_3_12),
    .valid_o_gather_pe              (gather_valid_o_3_12),
    .data_o_gather_pe               (gather_data_o_3_12),
    .ready_i_gather_pe              (gather_ready_i_3_12),

    .credit_upd                     (credit_upd[3][12])
);


network_interface #(
    .cast_out                       (cast_out_3_13),
    .gather_out                     (gather_out_3_13),
    .cast_sid                       (cast_sid_3_13),
    .gather_sid                     (gather_sid_3_13)
)ni_3_13(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[3][13]),
    .data_i_cast_nw                 (data_o_cast_nw[3][13]),
    .ready_o_cast_nw                (ready_i_cast_nw[3][13]),
    .valid_o_cast_nw                (valid_i_cast_nw[3][13]),
    .data_o_cast_nw                 (data_i_cast_nw[3][13]),
    .ready_i_cast_nw                (ready_o_cast_nw[3][13]),

    .valid_i_gather_nw              (valid_o_gather_nw[3][13]),
    .data_i_gather_nw               (data_o_gather_nw[3][13]),
    .ready_o_gather_nw              (ready_i_gather_nw[3][13]),
    .valid_o_gather_nw              (valid_i_gather_nw[3][13]),
    .data_o_gather_nw               (data_i_gather_nw[3][13]),
    .ready_i_gather_nw              (ready_o_gather_nw[3][13]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[3][13]),
    .data_i_merge_nw                (data_o_merge_nw[3][13]),
    .ready_o_merge_nw               (ready_i_merge_nw[3][13]),
    .valid_o_merge_nw               (valid_i_merge_nw[3][13]),
    .data_o_merge_nw                (data_i_merge_nw[3][13]),
    .ready_i_merge_nw               (ready_o_merge_nw[3][13]),

    .valid_i_cast_pe                (cast_valid_i_3_13),
    .data_i_cast_pe                 (cast_data_i_3_13),
    .ready_o_cast_pe                (cast_ready_o_3_13),
    .valid_o_cast_pe                (cast_valid_o_3_13),
    .data_o_cast_pe                 (cast_data_o_3_13),
    .ready_i_cast_pe                (cast_ready_i_3_13),

    .valid_i_merge_pe               (merge_valid_i_3_13),
    .data_i_merge_pe                (merge_data_i_3_13),
    .ready_o_merge_pe               (merge_ready_o_3_13),
    .valid_o_merge_pe               (merge_valid_o_3_13),
    .data_o_merge_pe                (merge_data_o_3_13),
    .ready_i_merge_pe               (merge_ready_i_3_13),

    .valid_i_gather_pe              (gather_valid_i_3_13),
    .data_i_gather_pe               (gather_data_i_3_13),
    .ready_o_gather_pe              (gather_ready_o_3_13),
    .valid_o_gather_pe              (gather_valid_o_3_13),
    .data_o_gather_pe               (gather_data_o_3_13),
    .ready_i_gather_pe              (gather_ready_i_3_13),

    .credit_upd                     (credit_upd[3][13])
);


network_interface #(
    .cast_out                       (cast_out_3_14),
    .gather_out                     (gather_out_3_14),
    .cast_sid                       (cast_sid_3_14),
    .gather_sid                     (gather_sid_3_14)
)ni_3_14(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[3][14]),
    .data_i_cast_nw                 (data_o_cast_nw[3][14]),
    .ready_o_cast_nw                (ready_i_cast_nw[3][14]),
    .valid_o_cast_nw                (valid_i_cast_nw[3][14]),
    .data_o_cast_nw                 (data_i_cast_nw[3][14]),
    .ready_i_cast_nw                (ready_o_cast_nw[3][14]),

    .valid_i_gather_nw              (valid_o_gather_nw[3][14]),
    .data_i_gather_nw               (data_o_gather_nw[3][14]),
    .ready_o_gather_nw              (ready_i_gather_nw[3][14]),
    .valid_o_gather_nw              (valid_i_gather_nw[3][14]),
    .data_o_gather_nw               (data_i_gather_nw[3][14]),
    .ready_i_gather_nw              (ready_o_gather_nw[3][14]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[3][14]),
    .data_i_merge_nw                (data_o_merge_nw[3][14]),
    .ready_o_merge_nw               (ready_i_merge_nw[3][14]),
    .valid_o_merge_nw               (valid_i_merge_nw[3][14]),
    .data_o_merge_nw                (data_i_merge_nw[3][14]),
    .ready_i_merge_nw               (ready_o_merge_nw[3][14]),

    .valid_i_cast_pe                (cast_valid_i_3_14),
    .data_i_cast_pe                 (cast_data_i_3_14),
    .ready_o_cast_pe                (cast_ready_o_3_14),
    .valid_o_cast_pe                (cast_valid_o_3_14),
    .data_o_cast_pe                 (cast_data_o_3_14),
    .ready_i_cast_pe                (cast_ready_i_3_14),

    .valid_i_merge_pe               (merge_valid_i_3_14),
    .data_i_merge_pe                (merge_data_i_3_14),
    .ready_o_merge_pe               (merge_ready_o_3_14),
    .valid_o_merge_pe               (merge_valid_o_3_14),
    .data_o_merge_pe                (merge_data_o_3_14),
    .ready_i_merge_pe               (merge_ready_i_3_14),

    .valid_i_gather_pe              (gather_valid_i_3_14),
    .data_i_gather_pe               (gather_data_i_3_14),
    .ready_o_gather_pe              (gather_ready_o_3_14),
    .valid_o_gather_pe              (gather_valid_o_3_14),
    .data_o_gather_pe               (gather_data_o_3_14),
    .ready_i_gather_pe              (gather_ready_i_3_14),

    .credit_upd                     (credit_upd[3][14])
);


network_interface #(
    .cast_out                       (cast_out_3_15),
    .gather_out                     (gather_out_3_15),
    .cast_sid                       (cast_sid_3_15),
    .gather_sid                     (gather_sid_3_15)
)ni_3_15(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[3][15]),
    .data_i_cast_nw                 (data_o_cast_nw[3][15]),
    .ready_o_cast_nw                (ready_i_cast_nw[3][15]),
    .valid_o_cast_nw                (valid_i_cast_nw[3][15]),
    .data_o_cast_nw                 (data_i_cast_nw[3][15]),
    .ready_i_cast_nw                (ready_o_cast_nw[3][15]),

    .valid_i_gather_nw              (valid_o_gather_nw[3][15]),
    .data_i_gather_nw               (data_o_gather_nw[3][15]),
    .ready_o_gather_nw              (ready_i_gather_nw[3][15]),
    .valid_o_gather_nw              (valid_i_gather_nw[3][15]),
    .data_o_gather_nw               (data_i_gather_nw[3][15]),
    .ready_i_gather_nw              (ready_o_gather_nw[3][15]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[3][15]),
    .data_i_merge_nw                (data_o_merge_nw[3][15]),
    .ready_o_merge_nw               (ready_i_merge_nw[3][15]),
    .valid_o_merge_nw               (valid_i_merge_nw[3][15]),
    .data_o_merge_nw                (data_i_merge_nw[3][15]),
    .ready_i_merge_nw               (ready_o_merge_nw[3][15]),

    .valid_i_cast_pe                (cast_valid_i_3_15),
    .data_i_cast_pe                 (cast_data_i_3_15),
    .ready_o_cast_pe                (cast_ready_o_3_15),
    .valid_o_cast_pe                (cast_valid_o_3_15),
    .data_o_cast_pe                 (cast_data_o_3_15),
    .ready_i_cast_pe                (cast_ready_i_3_15),

    .valid_i_merge_pe               (merge_valid_i_3_15),
    .data_i_merge_pe                (merge_data_i_3_15),
    .ready_o_merge_pe               (merge_ready_o_3_15),
    .valid_o_merge_pe               (merge_valid_o_3_15),
    .data_o_merge_pe                (merge_data_o_3_15),
    .ready_i_merge_pe               (merge_ready_i_3_15),

    .valid_i_gather_pe              (gather_valid_i_3_15),
    .data_i_gather_pe               (gather_data_i_3_15),
    .ready_o_gather_pe              (gather_ready_o_3_15),
    .valid_o_gather_pe              (gather_valid_o_3_15),
    .data_o_gather_pe               (gather_data_o_3_15),
    .ready_i_gather_pe              (gather_ready_i_3_15),

    .credit_upd                     (credit_upd[3][15])
);


network_interface #(
    .cast_out                       (cast_out_3_16),
    .gather_out                     (gather_out_3_16),
    .cast_sid                       (cast_sid_3_16),
    .gather_sid                     (gather_sid_3_16)
)ni_3_16(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[3][16]),
    .data_i_cast_nw                 (data_o_cast_nw[3][16]),
    .ready_o_cast_nw                (ready_i_cast_nw[3][16]),
    .valid_o_cast_nw                (valid_i_cast_nw[3][16]),
    .data_o_cast_nw                 (data_i_cast_nw[3][16]),
    .ready_i_cast_nw                (ready_o_cast_nw[3][16]),

    .valid_i_gather_nw              (valid_o_gather_nw[3][16]),
    .data_i_gather_nw               (data_o_gather_nw[3][16]),
    .ready_o_gather_nw              (ready_i_gather_nw[3][16]),
    .valid_o_gather_nw              (valid_i_gather_nw[3][16]),
    .data_o_gather_nw               (data_i_gather_nw[3][16]),
    .ready_i_gather_nw              (ready_o_gather_nw[3][16]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[3][16]),
    .data_i_merge_nw                (data_o_merge_nw[3][16]),
    .ready_o_merge_nw               (ready_i_merge_nw[3][16]),
    .valid_o_merge_nw               (valid_i_merge_nw[3][16]),
    .data_o_merge_nw                (data_i_merge_nw[3][16]),
    .ready_i_merge_nw               (ready_o_merge_nw[3][16]),

    .valid_i_cast_pe                (cast_valid_i_3_16),
    .data_i_cast_pe                 (cast_data_i_3_16),
    .ready_o_cast_pe                (cast_ready_o_3_16),
    .valid_o_cast_pe                (cast_valid_o_3_16),
    .data_o_cast_pe                 (cast_data_o_3_16),
    .ready_i_cast_pe                (cast_ready_i_3_16),

    .valid_i_merge_pe               (merge_valid_i_3_16),
    .data_i_merge_pe                (merge_data_i_3_16),
    .ready_o_merge_pe               (merge_ready_o_3_16),
    .valid_o_merge_pe               (merge_valid_o_3_16),
    .data_o_merge_pe                (merge_data_o_3_16),
    .ready_i_merge_pe               (merge_ready_i_3_16),

    .valid_i_gather_pe              (gather_valid_i_3_16),
    .data_i_gather_pe               (gather_data_i_3_16),
    .ready_o_gather_pe              (gather_ready_o_3_16),
    .valid_o_gather_pe              (gather_valid_o_3_16),
    .data_o_gather_pe               (gather_data_o_3_16),
    .ready_i_gather_pe              (gather_ready_i_3_16),

    .credit_upd                     (credit_upd[3][16])
);


network_interface #(
    .cast_out                       (cast_out_3_17),
    .gather_out                     (gather_out_3_17),
    .cast_sid                       (cast_sid_3_17),
    .gather_sid                     (gather_sid_3_17)
)ni_3_17(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[3][17]),
    .data_i_cast_nw                 (data_o_cast_nw[3][17]),
    .ready_o_cast_nw                (ready_i_cast_nw[3][17]),
    .valid_o_cast_nw                (valid_i_cast_nw[3][17]),
    .data_o_cast_nw                 (data_i_cast_nw[3][17]),
    .ready_i_cast_nw                (ready_o_cast_nw[3][17]),

    .valid_i_gather_nw              (valid_o_gather_nw[3][17]),
    .data_i_gather_nw               (data_o_gather_nw[3][17]),
    .ready_o_gather_nw              (ready_i_gather_nw[3][17]),
    .valid_o_gather_nw              (valid_i_gather_nw[3][17]),
    .data_o_gather_nw               (data_i_gather_nw[3][17]),
    .ready_i_gather_nw              (ready_o_gather_nw[3][17]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[3][17]),
    .data_i_merge_nw                (data_o_merge_nw[3][17]),
    .ready_o_merge_nw               (ready_i_merge_nw[3][17]),
    .valid_o_merge_nw               (valid_i_merge_nw[3][17]),
    .data_o_merge_nw                (data_i_merge_nw[3][17]),
    .ready_i_merge_nw               (ready_o_merge_nw[3][17]),

    .valid_i_cast_pe                (cast_valid_i_3_17),
    .data_i_cast_pe                 (cast_data_i_3_17),
    .ready_o_cast_pe                (cast_ready_o_3_17),
    .valid_o_cast_pe                (cast_valid_o_3_17),
    .data_o_cast_pe                 (cast_data_o_3_17),
    .ready_i_cast_pe                (cast_ready_i_3_17),

    .valid_i_merge_pe               (merge_valid_i_3_17),
    .data_i_merge_pe                (merge_data_i_3_17),
    .ready_o_merge_pe               (merge_ready_o_3_17),
    .valid_o_merge_pe               (merge_valid_o_3_17),
    .data_o_merge_pe                (merge_data_o_3_17),
    .ready_i_merge_pe               (merge_ready_i_3_17),

    .valid_i_gather_pe              (gather_valid_i_3_17),
    .data_i_gather_pe               (gather_data_i_3_17),
    .ready_o_gather_pe              (gather_ready_o_3_17),
    .valid_o_gather_pe              (gather_valid_o_3_17),
    .data_o_gather_pe               (gather_data_o_3_17),
    .ready_i_gather_pe              (gather_ready_i_3_17),

    .credit_upd                     (credit_upd[3][17])
);


network_interface #(
    .cast_out                       (cast_out_3_18),
    .gather_out                     (gather_out_3_18),
    .cast_sid                       (cast_sid_3_18),
    .gather_sid                     (gather_sid_3_18)
)ni_3_18(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[3][18]),
    .data_i_cast_nw                 (data_o_cast_nw[3][18]),
    .ready_o_cast_nw                (ready_i_cast_nw[3][18]),
    .valid_o_cast_nw                (valid_i_cast_nw[3][18]),
    .data_o_cast_nw                 (data_i_cast_nw[3][18]),
    .ready_i_cast_nw                (ready_o_cast_nw[3][18]),

    .valid_i_gather_nw              (valid_o_gather_nw[3][18]),
    .data_i_gather_nw               (data_o_gather_nw[3][18]),
    .ready_o_gather_nw              (ready_i_gather_nw[3][18]),
    .valid_o_gather_nw              (valid_i_gather_nw[3][18]),
    .data_o_gather_nw               (data_i_gather_nw[3][18]),
    .ready_i_gather_nw              (ready_o_gather_nw[3][18]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[3][18]),
    .data_i_merge_nw                (data_o_merge_nw[3][18]),
    .ready_o_merge_nw               (ready_i_merge_nw[3][18]),
    .valid_o_merge_nw               (valid_i_merge_nw[3][18]),
    .data_o_merge_nw                (data_i_merge_nw[3][18]),
    .ready_i_merge_nw               (ready_o_merge_nw[3][18]),

    .valid_i_cast_pe                (cast_valid_i_3_18),
    .data_i_cast_pe                 (cast_data_i_3_18),
    .ready_o_cast_pe                (cast_ready_o_3_18),
    .valid_o_cast_pe                (cast_valid_o_3_18),
    .data_o_cast_pe                 (cast_data_o_3_18),
    .ready_i_cast_pe                (cast_ready_i_3_18),

    .valid_i_merge_pe               (merge_valid_i_3_18),
    .data_i_merge_pe                (merge_data_i_3_18),
    .ready_o_merge_pe               (merge_ready_o_3_18),
    .valid_o_merge_pe               (merge_valid_o_3_18),
    .data_o_merge_pe                (merge_data_o_3_18),
    .ready_i_merge_pe               (merge_ready_i_3_18),

    .valid_i_gather_pe              (gather_valid_i_3_18),
    .data_i_gather_pe               (gather_data_i_3_18),
    .ready_o_gather_pe              (gather_ready_o_3_18),
    .valid_o_gather_pe              (gather_valid_o_3_18),
    .data_o_gather_pe               (gather_data_o_3_18),
    .ready_i_gather_pe              (gather_ready_i_3_18),

    .credit_upd                     (credit_upd[3][18])
);


network_interface #(
    .cast_out                       (cast_out_3_19),
    .gather_out                     (gather_out_3_19),
    .cast_sid                       (cast_sid_3_19),
    .gather_sid                     (gather_sid_3_19)
)ni_3_19(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[3][19]),
    .data_i_cast_nw                 (data_o_cast_nw[3][19]),
    .ready_o_cast_nw                (ready_i_cast_nw[3][19]),
    .valid_o_cast_nw                (valid_i_cast_nw[3][19]),
    .data_o_cast_nw                 (data_i_cast_nw[3][19]),
    .ready_i_cast_nw                (ready_o_cast_nw[3][19]),

    .valid_i_gather_nw              (valid_o_gather_nw[3][19]),
    .data_i_gather_nw               (data_o_gather_nw[3][19]),
    .ready_o_gather_nw              (ready_i_gather_nw[3][19]),
    .valid_o_gather_nw              (valid_i_gather_nw[3][19]),
    .data_o_gather_nw               (data_i_gather_nw[3][19]),
    .ready_i_gather_nw              (ready_o_gather_nw[3][19]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[3][19]),
    .data_i_merge_nw                (data_o_merge_nw[3][19]),
    .ready_o_merge_nw               (ready_i_merge_nw[3][19]),
    .valid_o_merge_nw               (valid_i_merge_nw[3][19]),
    .data_o_merge_nw                (data_i_merge_nw[3][19]),
    .ready_i_merge_nw               (ready_o_merge_nw[3][19]),

    .valid_i_cast_pe                (cast_valid_i_3_19),
    .data_i_cast_pe                 (cast_data_i_3_19),
    .ready_o_cast_pe                (cast_ready_o_3_19),
    .valid_o_cast_pe                (cast_valid_o_3_19),
    .data_o_cast_pe                 (cast_data_o_3_19),
    .ready_i_cast_pe                (cast_ready_i_3_19),

    .valid_i_merge_pe               (merge_valid_i_3_19),
    .data_i_merge_pe                (merge_data_i_3_19),
    .ready_o_merge_pe               (merge_ready_o_3_19),
    .valid_o_merge_pe               (merge_valid_o_3_19),
    .data_o_merge_pe                (merge_data_o_3_19),
    .ready_i_merge_pe               (merge_ready_i_3_19),

    .valid_i_gather_pe              (gather_valid_i_3_19),
    .data_i_gather_pe               (gather_data_i_3_19),
    .ready_o_gather_pe              (gather_ready_o_3_19),
    .valid_o_gather_pe              (gather_valid_o_3_19),
    .data_o_gather_pe               (gather_data_o_3_19),
    .ready_i_gather_pe              (gather_ready_i_3_19),

    .credit_upd                     (credit_upd[3][19])
);


network_interface #(
    .cast_out                       (cast_out_3_20),
    .gather_out                     (gather_out_3_20),
    .cast_sid                       (cast_sid_3_20),
    .gather_sid                     (gather_sid_3_20)
)ni_3_20(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[3][20]),
    .data_i_cast_nw                 (data_o_cast_nw[3][20]),
    .ready_o_cast_nw                (ready_i_cast_nw[3][20]),
    .valid_o_cast_nw                (valid_i_cast_nw[3][20]),
    .data_o_cast_nw                 (data_i_cast_nw[3][20]),
    .ready_i_cast_nw                (ready_o_cast_nw[3][20]),

    .valid_i_gather_nw              (valid_o_gather_nw[3][20]),
    .data_i_gather_nw               (data_o_gather_nw[3][20]),
    .ready_o_gather_nw              (ready_i_gather_nw[3][20]),
    .valid_o_gather_nw              (valid_i_gather_nw[3][20]),
    .data_o_gather_nw               (data_i_gather_nw[3][20]),
    .ready_i_gather_nw              (ready_o_gather_nw[3][20]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[3][20]),
    .data_i_merge_nw                (data_o_merge_nw[3][20]),
    .ready_o_merge_nw               (ready_i_merge_nw[3][20]),
    .valid_o_merge_nw               (valid_i_merge_nw[3][20]),
    .data_o_merge_nw                (data_i_merge_nw[3][20]),
    .ready_i_merge_nw               (ready_o_merge_nw[3][20]),

    .valid_i_cast_pe                (cast_valid_i_3_20),
    .data_i_cast_pe                 (cast_data_i_3_20),
    .ready_o_cast_pe                (cast_ready_o_3_20),
    .valid_o_cast_pe                (cast_valid_o_3_20),
    .data_o_cast_pe                 (cast_data_o_3_20),
    .ready_i_cast_pe                (cast_ready_i_3_20),

    .valid_i_merge_pe               (merge_valid_i_3_20),
    .data_i_merge_pe                (merge_data_i_3_20),
    .ready_o_merge_pe               (merge_ready_o_3_20),
    .valid_o_merge_pe               (merge_valid_o_3_20),
    .data_o_merge_pe                (merge_data_o_3_20),
    .ready_i_merge_pe               (merge_ready_i_3_20),

    .valid_i_gather_pe              (gather_valid_i_3_20),
    .data_i_gather_pe               (gather_data_i_3_20),
    .ready_o_gather_pe              (gather_ready_o_3_20),
    .valid_o_gather_pe              (gather_valid_o_3_20),
    .data_o_gather_pe               (gather_data_o_3_20),
    .ready_i_gather_pe              (gather_ready_i_3_20),

    .credit_upd                     (credit_upd[3][20])
);


network_interface #(
    .cast_out                       (cast_out_3_21),
    .gather_out                     (gather_out_3_21),
    .cast_sid                       (cast_sid_3_21),
    .gather_sid                     (gather_sid_3_21)
)ni_3_21(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[3][21]),
    .data_i_cast_nw                 (data_o_cast_nw[3][21]),
    .ready_o_cast_nw                (ready_i_cast_nw[3][21]),
    .valid_o_cast_nw                (valid_i_cast_nw[3][21]),
    .data_o_cast_nw                 (data_i_cast_nw[3][21]),
    .ready_i_cast_nw                (ready_o_cast_nw[3][21]),

    .valid_i_gather_nw              (valid_o_gather_nw[3][21]),
    .data_i_gather_nw               (data_o_gather_nw[3][21]),
    .ready_o_gather_nw              (ready_i_gather_nw[3][21]),
    .valid_o_gather_nw              (valid_i_gather_nw[3][21]),
    .data_o_gather_nw               (data_i_gather_nw[3][21]),
    .ready_i_gather_nw              (ready_o_gather_nw[3][21]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[3][21]),
    .data_i_merge_nw                (data_o_merge_nw[3][21]),
    .ready_o_merge_nw               (ready_i_merge_nw[3][21]),
    .valid_o_merge_nw               (valid_i_merge_nw[3][21]),
    .data_o_merge_nw                (data_i_merge_nw[3][21]),
    .ready_i_merge_nw               (ready_o_merge_nw[3][21]),

    .valid_i_cast_pe                (cast_valid_i_3_21),
    .data_i_cast_pe                 (cast_data_i_3_21),
    .ready_o_cast_pe                (cast_ready_o_3_21),
    .valid_o_cast_pe                (cast_valid_o_3_21),
    .data_o_cast_pe                 (cast_data_o_3_21),
    .ready_i_cast_pe                (cast_ready_i_3_21),

    .valid_i_merge_pe               (merge_valid_i_3_21),
    .data_i_merge_pe                (merge_data_i_3_21),
    .ready_o_merge_pe               (merge_ready_o_3_21),
    .valid_o_merge_pe               (merge_valid_o_3_21),
    .data_o_merge_pe                (merge_data_o_3_21),
    .ready_i_merge_pe               (merge_ready_i_3_21),

    .valid_i_gather_pe              (gather_valid_i_3_21),
    .data_i_gather_pe               (gather_data_i_3_21),
    .ready_o_gather_pe              (gather_ready_o_3_21),
    .valid_o_gather_pe              (gather_valid_o_3_21),
    .data_o_gather_pe               (gather_data_o_3_21),
    .ready_i_gather_pe              (gather_ready_i_3_21),

    .credit_upd                     (credit_upd[3][21])
);


network_interface #(
    .cast_out                       (cast_out_3_22),
    .gather_out                     (gather_out_3_22),
    .cast_sid                       (cast_sid_3_22),
    .gather_sid                     (gather_sid_3_22)
)ni_3_22(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[3][22]),
    .data_i_cast_nw                 (data_o_cast_nw[3][22]),
    .ready_o_cast_nw                (ready_i_cast_nw[3][22]),
    .valid_o_cast_nw                (valid_i_cast_nw[3][22]),
    .data_o_cast_nw                 (data_i_cast_nw[3][22]),
    .ready_i_cast_nw                (ready_o_cast_nw[3][22]),

    .valid_i_gather_nw              (valid_o_gather_nw[3][22]),
    .data_i_gather_nw               (data_o_gather_nw[3][22]),
    .ready_o_gather_nw              (ready_i_gather_nw[3][22]),
    .valid_o_gather_nw              (valid_i_gather_nw[3][22]),
    .data_o_gather_nw               (data_i_gather_nw[3][22]),
    .ready_i_gather_nw              (ready_o_gather_nw[3][22]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[3][22]),
    .data_i_merge_nw                (data_o_merge_nw[3][22]),
    .ready_o_merge_nw               (ready_i_merge_nw[3][22]),
    .valid_o_merge_nw               (valid_i_merge_nw[3][22]),
    .data_o_merge_nw                (data_i_merge_nw[3][22]),
    .ready_i_merge_nw               (ready_o_merge_nw[3][22]),

    .valid_i_cast_pe                (cast_valid_i_3_22),
    .data_i_cast_pe                 (cast_data_i_3_22),
    .ready_o_cast_pe                (cast_ready_o_3_22),
    .valid_o_cast_pe                (cast_valid_o_3_22),
    .data_o_cast_pe                 (cast_data_o_3_22),
    .ready_i_cast_pe                (cast_ready_i_3_22),

    .valid_i_merge_pe               (merge_valid_i_3_22),
    .data_i_merge_pe                (merge_data_i_3_22),
    .ready_o_merge_pe               (merge_ready_o_3_22),
    .valid_o_merge_pe               (merge_valid_o_3_22),
    .data_o_merge_pe                (merge_data_o_3_22),
    .ready_i_merge_pe               (merge_ready_i_3_22),

    .valid_i_gather_pe              (gather_valid_i_3_22),
    .data_i_gather_pe               (gather_data_i_3_22),
    .ready_o_gather_pe              (gather_ready_o_3_22),
    .valid_o_gather_pe              (gather_valid_o_3_22),
    .data_o_gather_pe               (gather_data_o_3_22),
    .ready_i_gather_pe              (gather_ready_i_3_22),

    .credit_upd                     (credit_upd[3][22])
);


network_interface #(
    .cast_out                       (cast_out_3_23),
    .gather_out                     (gather_out_3_23),
    .cast_sid                       (cast_sid_3_23),
    .gather_sid                     (gather_sid_3_23)
)ni_3_23(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[3][23]),
    .data_i_cast_nw                 (data_o_cast_nw[3][23]),
    .ready_o_cast_nw                (ready_i_cast_nw[3][23]),
    .valid_o_cast_nw                (valid_i_cast_nw[3][23]),
    .data_o_cast_nw                 (data_i_cast_nw[3][23]),
    .ready_i_cast_nw                (ready_o_cast_nw[3][23]),

    .valid_i_gather_nw              (valid_o_gather_nw[3][23]),
    .data_i_gather_nw               (data_o_gather_nw[3][23]),
    .ready_o_gather_nw              (ready_i_gather_nw[3][23]),
    .valid_o_gather_nw              (valid_i_gather_nw[3][23]),
    .data_o_gather_nw               (data_i_gather_nw[3][23]),
    .ready_i_gather_nw              (ready_o_gather_nw[3][23]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[3][23]),
    .data_i_merge_nw                (data_o_merge_nw[3][23]),
    .ready_o_merge_nw               (ready_i_merge_nw[3][23]),
    .valid_o_merge_nw               (valid_i_merge_nw[3][23]),
    .data_o_merge_nw                (data_i_merge_nw[3][23]),
    .ready_i_merge_nw               (ready_o_merge_nw[3][23]),

    .valid_i_cast_pe                (cast_valid_i_3_23),
    .data_i_cast_pe                 (cast_data_i_3_23),
    .ready_o_cast_pe                (cast_ready_o_3_23),
    .valid_o_cast_pe                (cast_valid_o_3_23),
    .data_o_cast_pe                 (cast_data_o_3_23),
    .ready_i_cast_pe                (cast_ready_i_3_23),

    .valid_i_merge_pe               (merge_valid_i_3_23),
    .data_i_merge_pe                (merge_data_i_3_23),
    .ready_o_merge_pe               (merge_ready_o_3_23),
    .valid_o_merge_pe               (merge_valid_o_3_23),
    .data_o_merge_pe                (merge_data_o_3_23),
    .ready_i_merge_pe               (merge_ready_i_3_23),

    .valid_i_gather_pe              (gather_valid_i_3_23),
    .data_i_gather_pe               (gather_data_i_3_23),
    .ready_o_gather_pe              (gather_ready_o_3_23),
    .valid_o_gather_pe              (gather_valid_o_3_23),
    .data_o_gather_pe               (gather_data_o_3_23),
    .ready_i_gather_pe              (gather_ready_i_3_23),

    .credit_upd                     (credit_upd[3][23])
);


network_interface #(
    .cast_out                       (cast_out_3_24),
    .gather_out                     (gather_out_3_24),
    .cast_sid                       (cast_sid_3_24),
    .gather_sid                     (gather_sid_3_24)
)ni_3_24(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[3][24]),
    .data_i_cast_nw                 (data_o_cast_nw[3][24]),
    .ready_o_cast_nw                (ready_i_cast_nw[3][24]),
    .valid_o_cast_nw                (valid_i_cast_nw[3][24]),
    .data_o_cast_nw                 (data_i_cast_nw[3][24]),
    .ready_i_cast_nw                (ready_o_cast_nw[3][24]),

    .valid_i_gather_nw              (valid_o_gather_nw[3][24]),
    .data_i_gather_nw               (data_o_gather_nw[3][24]),
    .ready_o_gather_nw              (ready_i_gather_nw[3][24]),
    .valid_o_gather_nw              (valid_i_gather_nw[3][24]),
    .data_o_gather_nw               (data_i_gather_nw[3][24]),
    .ready_i_gather_nw              (ready_o_gather_nw[3][24]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[3][24]),
    .data_i_merge_nw                (data_o_merge_nw[3][24]),
    .ready_o_merge_nw               (ready_i_merge_nw[3][24]),
    .valid_o_merge_nw               (valid_i_merge_nw[3][24]),
    .data_o_merge_nw                (data_i_merge_nw[3][24]),
    .ready_i_merge_nw               (ready_o_merge_nw[3][24]),

    .valid_i_cast_pe                (cast_valid_i_3_24),
    .data_i_cast_pe                 (cast_data_i_3_24),
    .ready_o_cast_pe                (cast_ready_o_3_24),
    .valid_o_cast_pe                (cast_valid_o_3_24),
    .data_o_cast_pe                 (cast_data_o_3_24),
    .ready_i_cast_pe                (cast_ready_i_3_24),

    .valid_i_merge_pe               (merge_valid_i_3_24),
    .data_i_merge_pe                (merge_data_i_3_24),
    .ready_o_merge_pe               (merge_ready_o_3_24),
    .valid_o_merge_pe               (merge_valid_o_3_24),
    .data_o_merge_pe                (merge_data_o_3_24),
    .ready_i_merge_pe               (merge_ready_i_3_24),

    .valid_i_gather_pe              (gather_valid_i_3_24),
    .data_i_gather_pe               (gather_data_i_3_24),
    .ready_o_gather_pe              (gather_ready_o_3_24),
    .valid_o_gather_pe              (gather_valid_o_3_24),
    .data_o_gather_pe               (gather_data_o_3_24),
    .ready_i_gather_pe              (gather_ready_i_3_24),

    .credit_upd                     (credit_upd[3][24])
);


network_interface #(
    .cast_out                       (cast_out_4_0),
    .gather_out                     (gather_out_4_0),
    .cast_sid                       (cast_sid_4_0),
    .gather_sid                     (gather_sid_4_0)
)ni_4_0(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[4][0]),
    .data_i_cast_nw                 (data_o_cast_nw[4][0]),
    .ready_o_cast_nw                (ready_i_cast_nw[4][0]),
    .valid_o_cast_nw                (valid_i_cast_nw[4][0]),
    .data_o_cast_nw                 (data_i_cast_nw[4][0]),
    .ready_i_cast_nw                (ready_o_cast_nw[4][0]),

    .valid_i_gather_nw              (valid_o_gather_nw[4][0]),
    .data_i_gather_nw               (data_o_gather_nw[4][0]),
    .ready_o_gather_nw              (ready_i_gather_nw[4][0]),
    .valid_o_gather_nw              (valid_i_gather_nw[4][0]),
    .data_o_gather_nw               (data_i_gather_nw[4][0]),
    .ready_i_gather_nw              (ready_o_gather_nw[4][0]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[4][0]),
    .data_i_merge_nw                (data_o_merge_nw[4][0]),
    .ready_o_merge_nw               (ready_i_merge_nw[4][0]),
    .valid_o_merge_nw               (valid_i_merge_nw[4][0]),
    .data_o_merge_nw                (data_i_merge_nw[4][0]),
    .ready_i_merge_nw               (ready_o_merge_nw[4][0]),

    .valid_i_cast_pe                (cast_valid_i_4_0),
    .data_i_cast_pe                 (cast_data_i_4_0),
    .ready_o_cast_pe                (cast_ready_o_4_0),
    .valid_o_cast_pe                (cast_valid_o_4_0),
    .data_o_cast_pe                 (cast_data_o_4_0),
    .ready_i_cast_pe                (cast_ready_i_4_0),

    .valid_i_merge_pe               (merge_valid_i_4_0),
    .data_i_merge_pe                (merge_data_i_4_0),
    .ready_o_merge_pe               (merge_ready_o_4_0),
    .valid_o_merge_pe               (merge_valid_o_4_0),
    .data_o_merge_pe                (merge_data_o_4_0),
    .ready_i_merge_pe               (merge_ready_i_4_0),

    .valid_i_gather_pe              (gather_valid_i_4_0),
    .data_i_gather_pe               (gather_data_i_4_0),
    .ready_o_gather_pe              (gather_ready_o_4_0),
    .valid_o_gather_pe              (gather_valid_o_4_0),
    .data_o_gather_pe               (gather_data_o_4_0),
    .ready_i_gather_pe              (gather_ready_i_4_0),

    .credit_upd                     (credit_upd[4][0])
);


network_interface #(
    .cast_out                       (cast_out_4_1),
    .gather_out                     (gather_out_4_1),
    .cast_sid                       (cast_sid_4_1),
    .gather_sid                     (gather_sid_4_1)
)ni_4_1(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[4][1]),
    .data_i_cast_nw                 (data_o_cast_nw[4][1]),
    .ready_o_cast_nw                (ready_i_cast_nw[4][1]),
    .valid_o_cast_nw                (valid_i_cast_nw[4][1]),
    .data_o_cast_nw                 (data_i_cast_nw[4][1]),
    .ready_i_cast_nw                (ready_o_cast_nw[4][1]),

    .valid_i_gather_nw              (valid_o_gather_nw[4][1]),
    .data_i_gather_nw               (data_o_gather_nw[4][1]),
    .ready_o_gather_nw              (ready_i_gather_nw[4][1]),
    .valid_o_gather_nw              (valid_i_gather_nw[4][1]),
    .data_o_gather_nw               (data_i_gather_nw[4][1]),
    .ready_i_gather_nw              (ready_o_gather_nw[4][1]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[4][1]),
    .data_i_merge_nw                (data_o_merge_nw[4][1]),
    .ready_o_merge_nw               (ready_i_merge_nw[4][1]),
    .valid_o_merge_nw               (valid_i_merge_nw[4][1]),
    .data_o_merge_nw                (data_i_merge_nw[4][1]),
    .ready_i_merge_nw               (ready_o_merge_nw[4][1]),

    .valid_i_cast_pe                (cast_valid_i_4_1),
    .data_i_cast_pe                 (cast_data_i_4_1),
    .ready_o_cast_pe                (cast_ready_o_4_1),
    .valid_o_cast_pe                (cast_valid_o_4_1),
    .data_o_cast_pe                 (cast_data_o_4_1),
    .ready_i_cast_pe                (cast_ready_i_4_1),

    .valid_i_merge_pe               (merge_valid_i_4_1),
    .data_i_merge_pe                (merge_data_i_4_1),
    .ready_o_merge_pe               (merge_ready_o_4_1),
    .valid_o_merge_pe               (merge_valid_o_4_1),
    .data_o_merge_pe                (merge_data_o_4_1),
    .ready_i_merge_pe               (merge_ready_i_4_1),

    .valid_i_gather_pe              (gather_valid_i_4_1),
    .data_i_gather_pe               (gather_data_i_4_1),
    .ready_o_gather_pe              (gather_ready_o_4_1),
    .valid_o_gather_pe              (gather_valid_o_4_1),
    .data_o_gather_pe               (gather_data_o_4_1),
    .ready_i_gather_pe              (gather_ready_i_4_1),

    .credit_upd                     (credit_upd[4][1])
);


network_interface #(
    .cast_out                       (cast_out_4_2),
    .gather_out                     (gather_out_4_2),
    .cast_sid                       (cast_sid_4_2),
    .gather_sid                     (gather_sid_4_2)
)ni_4_2(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[4][2]),
    .data_i_cast_nw                 (data_o_cast_nw[4][2]),
    .ready_o_cast_nw                (ready_i_cast_nw[4][2]),
    .valid_o_cast_nw                (valid_i_cast_nw[4][2]),
    .data_o_cast_nw                 (data_i_cast_nw[4][2]),
    .ready_i_cast_nw                (ready_o_cast_nw[4][2]),

    .valid_i_gather_nw              (valid_o_gather_nw[4][2]),
    .data_i_gather_nw               (data_o_gather_nw[4][2]),
    .ready_o_gather_nw              (ready_i_gather_nw[4][2]),
    .valid_o_gather_nw              (valid_i_gather_nw[4][2]),
    .data_o_gather_nw               (data_i_gather_nw[4][2]),
    .ready_i_gather_nw              (ready_o_gather_nw[4][2]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[4][2]),
    .data_i_merge_nw                (data_o_merge_nw[4][2]),
    .ready_o_merge_nw               (ready_i_merge_nw[4][2]),
    .valid_o_merge_nw               (valid_i_merge_nw[4][2]),
    .data_o_merge_nw                (data_i_merge_nw[4][2]),
    .ready_i_merge_nw               (ready_o_merge_nw[4][2]),

    .valid_i_cast_pe                (cast_valid_i_4_2),
    .data_i_cast_pe                 (cast_data_i_4_2),
    .ready_o_cast_pe                (cast_ready_o_4_2),
    .valid_o_cast_pe                (cast_valid_o_4_2),
    .data_o_cast_pe                 (cast_data_o_4_2),
    .ready_i_cast_pe                (cast_ready_i_4_2),

    .valid_i_merge_pe               (merge_valid_i_4_2),
    .data_i_merge_pe                (merge_data_i_4_2),
    .ready_o_merge_pe               (merge_ready_o_4_2),
    .valid_o_merge_pe               (merge_valid_o_4_2),
    .data_o_merge_pe                (merge_data_o_4_2),
    .ready_i_merge_pe               (merge_ready_i_4_2),

    .valid_i_gather_pe              (gather_valid_i_4_2),
    .data_i_gather_pe               (gather_data_i_4_2),
    .ready_o_gather_pe              (gather_ready_o_4_2),
    .valid_o_gather_pe              (gather_valid_o_4_2),
    .data_o_gather_pe               (gather_data_o_4_2),
    .ready_i_gather_pe              (gather_ready_i_4_2),

    .credit_upd                     (credit_upd[4][2])
);


network_interface #(
    .cast_out                       (cast_out_4_3),
    .gather_out                     (gather_out_4_3),
    .cast_sid                       (cast_sid_4_3),
    .gather_sid                     (gather_sid_4_3)
)ni_4_3(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[4][3]),
    .data_i_cast_nw                 (data_o_cast_nw[4][3]),
    .ready_o_cast_nw                (ready_i_cast_nw[4][3]),
    .valid_o_cast_nw                (valid_i_cast_nw[4][3]),
    .data_o_cast_nw                 (data_i_cast_nw[4][3]),
    .ready_i_cast_nw                (ready_o_cast_nw[4][3]),

    .valid_i_gather_nw              (valid_o_gather_nw[4][3]),
    .data_i_gather_nw               (data_o_gather_nw[4][3]),
    .ready_o_gather_nw              (ready_i_gather_nw[4][3]),
    .valid_o_gather_nw              (valid_i_gather_nw[4][3]),
    .data_o_gather_nw               (data_i_gather_nw[4][3]),
    .ready_i_gather_nw              (ready_o_gather_nw[4][3]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[4][3]),
    .data_i_merge_nw                (data_o_merge_nw[4][3]),
    .ready_o_merge_nw               (ready_i_merge_nw[4][3]),
    .valid_o_merge_nw               (valid_i_merge_nw[4][3]),
    .data_o_merge_nw                (data_i_merge_nw[4][3]),
    .ready_i_merge_nw               (ready_o_merge_nw[4][3]),

    .valid_i_cast_pe                (cast_valid_i_4_3),
    .data_i_cast_pe                 (cast_data_i_4_3),
    .ready_o_cast_pe                (cast_ready_o_4_3),
    .valid_o_cast_pe                (cast_valid_o_4_3),
    .data_o_cast_pe                 (cast_data_o_4_3),
    .ready_i_cast_pe                (cast_ready_i_4_3),

    .valid_i_merge_pe               (merge_valid_i_4_3),
    .data_i_merge_pe                (merge_data_i_4_3),
    .ready_o_merge_pe               (merge_ready_o_4_3),
    .valid_o_merge_pe               (merge_valid_o_4_3),
    .data_o_merge_pe                (merge_data_o_4_3),
    .ready_i_merge_pe               (merge_ready_i_4_3),

    .valid_i_gather_pe              (gather_valid_i_4_3),
    .data_i_gather_pe               (gather_data_i_4_3),
    .ready_o_gather_pe              (gather_ready_o_4_3),
    .valid_o_gather_pe              (gather_valid_o_4_3),
    .data_o_gather_pe               (gather_data_o_4_3),
    .ready_i_gather_pe              (gather_ready_i_4_3),

    .credit_upd                     (credit_upd[4][3])
);


network_interface #(
    .cast_out                       (cast_out_4_4),
    .gather_out                     (gather_out_4_4),
    .cast_sid                       (cast_sid_4_4),
    .gather_sid                     (gather_sid_4_4)
)ni_4_4(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[4][4]),
    .data_i_cast_nw                 (data_o_cast_nw[4][4]),
    .ready_o_cast_nw                (ready_i_cast_nw[4][4]),
    .valid_o_cast_nw                (valid_i_cast_nw[4][4]),
    .data_o_cast_nw                 (data_i_cast_nw[4][4]),
    .ready_i_cast_nw                (ready_o_cast_nw[4][4]),

    .valid_i_gather_nw              (valid_o_gather_nw[4][4]),
    .data_i_gather_nw               (data_o_gather_nw[4][4]),
    .ready_o_gather_nw              (ready_i_gather_nw[4][4]),
    .valid_o_gather_nw              (valid_i_gather_nw[4][4]),
    .data_o_gather_nw               (data_i_gather_nw[4][4]),
    .ready_i_gather_nw              (ready_o_gather_nw[4][4]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[4][4]),
    .data_i_merge_nw                (data_o_merge_nw[4][4]),
    .ready_o_merge_nw               (ready_i_merge_nw[4][4]),
    .valid_o_merge_nw               (valid_i_merge_nw[4][4]),
    .data_o_merge_nw                (data_i_merge_nw[4][4]),
    .ready_i_merge_nw               (ready_o_merge_nw[4][4]),

    .valid_i_cast_pe                (cast_valid_i_4_4),
    .data_i_cast_pe                 (cast_data_i_4_4),
    .ready_o_cast_pe                (cast_ready_o_4_4),
    .valid_o_cast_pe                (cast_valid_o_4_4),
    .data_o_cast_pe                 (cast_data_o_4_4),
    .ready_i_cast_pe                (cast_ready_i_4_4),

    .valid_i_merge_pe               (merge_valid_i_4_4),
    .data_i_merge_pe                (merge_data_i_4_4),
    .ready_o_merge_pe               (merge_ready_o_4_4),
    .valid_o_merge_pe               (merge_valid_o_4_4),
    .data_o_merge_pe                (merge_data_o_4_4),
    .ready_i_merge_pe               (merge_ready_i_4_4),

    .valid_i_gather_pe              (gather_valid_i_4_4),
    .data_i_gather_pe               (gather_data_i_4_4),
    .ready_o_gather_pe              (gather_ready_o_4_4),
    .valid_o_gather_pe              (gather_valid_o_4_4),
    .data_o_gather_pe               (gather_data_o_4_4),
    .ready_i_gather_pe              (gather_ready_i_4_4),

    .credit_upd                     (credit_upd[4][4])
);


network_interface #(
    .cast_out                       (cast_out_4_5),
    .gather_out                     (gather_out_4_5),
    .cast_sid                       (cast_sid_4_5),
    .gather_sid                     (gather_sid_4_5)
)ni_4_5(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[4][5]),
    .data_i_cast_nw                 (data_o_cast_nw[4][5]),
    .ready_o_cast_nw                (ready_i_cast_nw[4][5]),
    .valid_o_cast_nw                (valid_i_cast_nw[4][5]),
    .data_o_cast_nw                 (data_i_cast_nw[4][5]),
    .ready_i_cast_nw                (ready_o_cast_nw[4][5]),

    .valid_i_gather_nw              (valid_o_gather_nw[4][5]),
    .data_i_gather_nw               (data_o_gather_nw[4][5]),
    .ready_o_gather_nw              (ready_i_gather_nw[4][5]),
    .valid_o_gather_nw              (valid_i_gather_nw[4][5]),
    .data_o_gather_nw               (data_i_gather_nw[4][5]),
    .ready_i_gather_nw              (ready_o_gather_nw[4][5]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[4][5]),
    .data_i_merge_nw                (data_o_merge_nw[4][5]),
    .ready_o_merge_nw               (ready_i_merge_nw[4][5]),
    .valid_o_merge_nw               (valid_i_merge_nw[4][5]),
    .data_o_merge_nw                (data_i_merge_nw[4][5]),
    .ready_i_merge_nw               (ready_o_merge_nw[4][5]),

    .valid_i_cast_pe                (cast_valid_i_4_5),
    .data_i_cast_pe                 (cast_data_i_4_5),
    .ready_o_cast_pe                (cast_ready_o_4_5),
    .valid_o_cast_pe                (cast_valid_o_4_5),
    .data_o_cast_pe                 (cast_data_o_4_5),
    .ready_i_cast_pe                (cast_ready_i_4_5),

    .valid_i_merge_pe               (merge_valid_i_4_5),
    .data_i_merge_pe                (merge_data_i_4_5),
    .ready_o_merge_pe               (merge_ready_o_4_5),
    .valid_o_merge_pe               (merge_valid_o_4_5),
    .data_o_merge_pe                (merge_data_o_4_5),
    .ready_i_merge_pe               (merge_ready_i_4_5),

    .valid_i_gather_pe              (gather_valid_i_4_5),
    .data_i_gather_pe               (gather_data_i_4_5),
    .ready_o_gather_pe              (gather_ready_o_4_5),
    .valid_o_gather_pe              (gather_valid_o_4_5),
    .data_o_gather_pe               (gather_data_o_4_5),
    .ready_i_gather_pe              (gather_ready_i_4_5),

    .credit_upd                     (credit_upd[4][5])
);


network_interface #(
    .cast_out                       (cast_out_4_6),
    .gather_out                     (gather_out_4_6),
    .cast_sid                       (cast_sid_4_6),
    .gather_sid                     (gather_sid_4_6)
)ni_4_6(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[4][6]),
    .data_i_cast_nw                 (data_o_cast_nw[4][6]),
    .ready_o_cast_nw                (ready_i_cast_nw[4][6]),
    .valid_o_cast_nw                (valid_i_cast_nw[4][6]),
    .data_o_cast_nw                 (data_i_cast_nw[4][6]),
    .ready_i_cast_nw                (ready_o_cast_nw[4][6]),

    .valid_i_gather_nw              (valid_o_gather_nw[4][6]),
    .data_i_gather_nw               (data_o_gather_nw[4][6]),
    .ready_o_gather_nw              (ready_i_gather_nw[4][6]),
    .valid_o_gather_nw              (valid_i_gather_nw[4][6]),
    .data_o_gather_nw               (data_i_gather_nw[4][6]),
    .ready_i_gather_nw              (ready_o_gather_nw[4][6]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[4][6]),
    .data_i_merge_nw                (data_o_merge_nw[4][6]),
    .ready_o_merge_nw               (ready_i_merge_nw[4][6]),
    .valid_o_merge_nw               (valid_i_merge_nw[4][6]),
    .data_o_merge_nw                (data_i_merge_nw[4][6]),
    .ready_i_merge_nw               (ready_o_merge_nw[4][6]),

    .valid_i_cast_pe                (cast_valid_i_4_6),
    .data_i_cast_pe                 (cast_data_i_4_6),
    .ready_o_cast_pe                (cast_ready_o_4_6),
    .valid_o_cast_pe                (cast_valid_o_4_6),
    .data_o_cast_pe                 (cast_data_o_4_6),
    .ready_i_cast_pe                (cast_ready_i_4_6),

    .valid_i_merge_pe               (merge_valid_i_4_6),
    .data_i_merge_pe                (merge_data_i_4_6),
    .ready_o_merge_pe               (merge_ready_o_4_6),
    .valid_o_merge_pe               (merge_valid_o_4_6),
    .data_o_merge_pe                (merge_data_o_4_6),
    .ready_i_merge_pe               (merge_ready_i_4_6),

    .valid_i_gather_pe              (gather_valid_i_4_6),
    .data_i_gather_pe               (gather_data_i_4_6),
    .ready_o_gather_pe              (gather_ready_o_4_6),
    .valid_o_gather_pe              (gather_valid_o_4_6),
    .data_o_gather_pe               (gather_data_o_4_6),
    .ready_i_gather_pe              (gather_ready_i_4_6),

    .credit_upd                     (credit_upd[4][6])
);


network_interface #(
    .cast_out                       (cast_out_4_7),
    .gather_out                     (gather_out_4_7),
    .cast_sid                       (cast_sid_4_7),
    .gather_sid                     (gather_sid_4_7)
)ni_4_7(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[4][7]),
    .data_i_cast_nw                 (data_o_cast_nw[4][7]),
    .ready_o_cast_nw                (ready_i_cast_nw[4][7]),
    .valid_o_cast_nw                (valid_i_cast_nw[4][7]),
    .data_o_cast_nw                 (data_i_cast_nw[4][7]),
    .ready_i_cast_nw                (ready_o_cast_nw[4][7]),

    .valid_i_gather_nw              (valid_o_gather_nw[4][7]),
    .data_i_gather_nw               (data_o_gather_nw[4][7]),
    .ready_o_gather_nw              (ready_i_gather_nw[4][7]),
    .valid_o_gather_nw              (valid_i_gather_nw[4][7]),
    .data_o_gather_nw               (data_i_gather_nw[4][7]),
    .ready_i_gather_nw              (ready_o_gather_nw[4][7]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[4][7]),
    .data_i_merge_nw                (data_o_merge_nw[4][7]),
    .ready_o_merge_nw               (ready_i_merge_nw[4][7]),
    .valid_o_merge_nw               (valid_i_merge_nw[4][7]),
    .data_o_merge_nw                (data_i_merge_nw[4][7]),
    .ready_i_merge_nw               (ready_o_merge_nw[4][7]),

    .valid_i_cast_pe                (cast_valid_i_4_7),
    .data_i_cast_pe                 (cast_data_i_4_7),
    .ready_o_cast_pe                (cast_ready_o_4_7),
    .valid_o_cast_pe                (cast_valid_o_4_7),
    .data_o_cast_pe                 (cast_data_o_4_7),
    .ready_i_cast_pe                (cast_ready_i_4_7),

    .valid_i_merge_pe               (merge_valid_i_4_7),
    .data_i_merge_pe                (merge_data_i_4_7),
    .ready_o_merge_pe               (merge_ready_o_4_7),
    .valid_o_merge_pe               (merge_valid_o_4_7),
    .data_o_merge_pe                (merge_data_o_4_7),
    .ready_i_merge_pe               (merge_ready_i_4_7),

    .valid_i_gather_pe              (gather_valid_i_4_7),
    .data_i_gather_pe               (gather_data_i_4_7),
    .ready_o_gather_pe              (gather_ready_o_4_7),
    .valid_o_gather_pe              (gather_valid_o_4_7),
    .data_o_gather_pe               (gather_data_o_4_7),
    .ready_i_gather_pe              (gather_ready_i_4_7),

    .credit_upd                     (credit_upd[4][7])
);


network_interface #(
    .cast_out                       (cast_out_4_8),
    .gather_out                     (gather_out_4_8),
    .cast_sid                       (cast_sid_4_8),
    .gather_sid                     (gather_sid_4_8)
)ni_4_8(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[4][8]),
    .data_i_cast_nw                 (data_o_cast_nw[4][8]),
    .ready_o_cast_nw                (ready_i_cast_nw[4][8]),
    .valid_o_cast_nw                (valid_i_cast_nw[4][8]),
    .data_o_cast_nw                 (data_i_cast_nw[4][8]),
    .ready_i_cast_nw                (ready_o_cast_nw[4][8]),

    .valid_i_gather_nw              (valid_o_gather_nw[4][8]),
    .data_i_gather_nw               (data_o_gather_nw[4][8]),
    .ready_o_gather_nw              (ready_i_gather_nw[4][8]),
    .valid_o_gather_nw              (valid_i_gather_nw[4][8]),
    .data_o_gather_nw               (data_i_gather_nw[4][8]),
    .ready_i_gather_nw              (ready_o_gather_nw[4][8]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[4][8]),
    .data_i_merge_nw                (data_o_merge_nw[4][8]),
    .ready_o_merge_nw               (ready_i_merge_nw[4][8]),
    .valid_o_merge_nw               (valid_i_merge_nw[4][8]),
    .data_o_merge_nw                (data_i_merge_nw[4][8]),
    .ready_i_merge_nw               (ready_o_merge_nw[4][8]),

    .valid_i_cast_pe                (cast_valid_i_4_8),
    .data_i_cast_pe                 (cast_data_i_4_8),
    .ready_o_cast_pe                (cast_ready_o_4_8),
    .valid_o_cast_pe                (cast_valid_o_4_8),
    .data_o_cast_pe                 (cast_data_o_4_8),
    .ready_i_cast_pe                (cast_ready_i_4_8),

    .valid_i_merge_pe               (merge_valid_i_4_8),
    .data_i_merge_pe                (merge_data_i_4_8),
    .ready_o_merge_pe               (merge_ready_o_4_8),
    .valid_o_merge_pe               (merge_valid_o_4_8),
    .data_o_merge_pe                (merge_data_o_4_8),
    .ready_i_merge_pe               (merge_ready_i_4_8),

    .valid_i_gather_pe              (gather_valid_i_4_8),
    .data_i_gather_pe               (gather_data_i_4_8),
    .ready_o_gather_pe              (gather_ready_o_4_8),
    .valid_o_gather_pe              (gather_valid_o_4_8),
    .data_o_gather_pe               (gather_data_o_4_8),
    .ready_i_gather_pe              (gather_ready_i_4_8),

    .credit_upd                     (credit_upd[4][8])
);


network_interface #(
    .cast_out                       (cast_out_4_9),
    .gather_out                     (gather_out_4_9),
    .cast_sid                       (cast_sid_4_9),
    .gather_sid                     (gather_sid_4_9)
)ni_4_9(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[4][9]),
    .data_i_cast_nw                 (data_o_cast_nw[4][9]),
    .ready_o_cast_nw                (ready_i_cast_nw[4][9]),
    .valid_o_cast_nw                (valid_i_cast_nw[4][9]),
    .data_o_cast_nw                 (data_i_cast_nw[4][9]),
    .ready_i_cast_nw                (ready_o_cast_nw[4][9]),

    .valid_i_gather_nw              (valid_o_gather_nw[4][9]),
    .data_i_gather_nw               (data_o_gather_nw[4][9]),
    .ready_o_gather_nw              (ready_i_gather_nw[4][9]),
    .valid_o_gather_nw              (valid_i_gather_nw[4][9]),
    .data_o_gather_nw               (data_i_gather_nw[4][9]),
    .ready_i_gather_nw              (ready_o_gather_nw[4][9]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[4][9]),
    .data_i_merge_nw                (data_o_merge_nw[4][9]),
    .ready_o_merge_nw               (ready_i_merge_nw[4][9]),
    .valid_o_merge_nw               (valid_i_merge_nw[4][9]),
    .data_o_merge_nw                (data_i_merge_nw[4][9]),
    .ready_i_merge_nw               (ready_o_merge_nw[4][9]),

    .valid_i_cast_pe                (cast_valid_i_4_9),
    .data_i_cast_pe                 (cast_data_i_4_9),
    .ready_o_cast_pe                (cast_ready_o_4_9),
    .valid_o_cast_pe                (cast_valid_o_4_9),
    .data_o_cast_pe                 (cast_data_o_4_9),
    .ready_i_cast_pe                (cast_ready_i_4_9),

    .valid_i_merge_pe               (merge_valid_i_4_9),
    .data_i_merge_pe                (merge_data_i_4_9),
    .ready_o_merge_pe               (merge_ready_o_4_9),
    .valid_o_merge_pe               (merge_valid_o_4_9),
    .data_o_merge_pe                (merge_data_o_4_9),
    .ready_i_merge_pe               (merge_ready_i_4_9),

    .valid_i_gather_pe              (gather_valid_i_4_9),
    .data_i_gather_pe               (gather_data_i_4_9),
    .ready_o_gather_pe              (gather_ready_o_4_9),
    .valid_o_gather_pe              (gather_valid_o_4_9),
    .data_o_gather_pe               (gather_data_o_4_9),
    .ready_i_gather_pe              (gather_ready_i_4_9),

    .credit_upd                     (credit_upd[4][9])
);


network_interface #(
    .cast_out                       (cast_out_4_10),
    .gather_out                     (gather_out_4_10),
    .cast_sid                       (cast_sid_4_10),
    .gather_sid                     (gather_sid_4_10)
)ni_4_10(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[4][10]),
    .data_i_cast_nw                 (data_o_cast_nw[4][10]),
    .ready_o_cast_nw                (ready_i_cast_nw[4][10]),
    .valid_o_cast_nw                (valid_i_cast_nw[4][10]),
    .data_o_cast_nw                 (data_i_cast_nw[4][10]),
    .ready_i_cast_nw                (ready_o_cast_nw[4][10]),

    .valid_i_gather_nw              (valid_o_gather_nw[4][10]),
    .data_i_gather_nw               (data_o_gather_nw[4][10]),
    .ready_o_gather_nw              (ready_i_gather_nw[4][10]),
    .valid_o_gather_nw              (valid_i_gather_nw[4][10]),
    .data_o_gather_nw               (data_i_gather_nw[4][10]),
    .ready_i_gather_nw              (ready_o_gather_nw[4][10]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[4][10]),
    .data_i_merge_nw                (data_o_merge_nw[4][10]),
    .ready_o_merge_nw               (ready_i_merge_nw[4][10]),
    .valid_o_merge_nw               (valid_i_merge_nw[4][10]),
    .data_o_merge_nw                (data_i_merge_nw[4][10]),
    .ready_i_merge_nw               (ready_o_merge_nw[4][10]),

    .valid_i_cast_pe                (cast_valid_i_4_10),
    .data_i_cast_pe                 (cast_data_i_4_10),
    .ready_o_cast_pe                (cast_ready_o_4_10),
    .valid_o_cast_pe                (cast_valid_o_4_10),
    .data_o_cast_pe                 (cast_data_o_4_10),
    .ready_i_cast_pe                (cast_ready_i_4_10),

    .valid_i_merge_pe               (merge_valid_i_4_10),
    .data_i_merge_pe                (merge_data_i_4_10),
    .ready_o_merge_pe               (merge_ready_o_4_10),
    .valid_o_merge_pe               (merge_valid_o_4_10),
    .data_o_merge_pe                (merge_data_o_4_10),
    .ready_i_merge_pe               (merge_ready_i_4_10),

    .valid_i_gather_pe              (gather_valid_i_4_10),
    .data_i_gather_pe               (gather_data_i_4_10),
    .ready_o_gather_pe              (gather_ready_o_4_10),
    .valid_o_gather_pe              (gather_valid_o_4_10),
    .data_o_gather_pe               (gather_data_o_4_10),
    .ready_i_gather_pe              (gather_ready_i_4_10),

    .credit_upd                     (credit_upd[4][10])
);


network_interface #(
    .cast_out                       (cast_out_4_11),
    .gather_out                     (gather_out_4_11),
    .cast_sid                       (cast_sid_4_11),
    .gather_sid                     (gather_sid_4_11)
)ni_4_11(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[4][11]),
    .data_i_cast_nw                 (data_o_cast_nw[4][11]),
    .ready_o_cast_nw                (ready_i_cast_nw[4][11]),
    .valid_o_cast_nw                (valid_i_cast_nw[4][11]),
    .data_o_cast_nw                 (data_i_cast_nw[4][11]),
    .ready_i_cast_nw                (ready_o_cast_nw[4][11]),

    .valid_i_gather_nw              (valid_o_gather_nw[4][11]),
    .data_i_gather_nw               (data_o_gather_nw[4][11]),
    .ready_o_gather_nw              (ready_i_gather_nw[4][11]),
    .valid_o_gather_nw              (valid_i_gather_nw[4][11]),
    .data_o_gather_nw               (data_i_gather_nw[4][11]),
    .ready_i_gather_nw              (ready_o_gather_nw[4][11]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[4][11]),
    .data_i_merge_nw                (data_o_merge_nw[4][11]),
    .ready_o_merge_nw               (ready_i_merge_nw[4][11]),
    .valid_o_merge_nw               (valid_i_merge_nw[4][11]),
    .data_o_merge_nw                (data_i_merge_nw[4][11]),
    .ready_i_merge_nw               (ready_o_merge_nw[4][11]),

    .valid_i_cast_pe                (cast_valid_i_4_11),
    .data_i_cast_pe                 (cast_data_i_4_11),
    .ready_o_cast_pe                (cast_ready_o_4_11),
    .valid_o_cast_pe                (cast_valid_o_4_11),
    .data_o_cast_pe                 (cast_data_o_4_11),
    .ready_i_cast_pe                (cast_ready_i_4_11),

    .valid_i_merge_pe               (merge_valid_i_4_11),
    .data_i_merge_pe                (merge_data_i_4_11),
    .ready_o_merge_pe               (merge_ready_o_4_11),
    .valid_o_merge_pe               (merge_valid_o_4_11),
    .data_o_merge_pe                (merge_data_o_4_11),
    .ready_i_merge_pe               (merge_ready_i_4_11),

    .valid_i_gather_pe              (gather_valid_i_4_11),
    .data_i_gather_pe               (gather_data_i_4_11),
    .ready_o_gather_pe              (gather_ready_o_4_11),
    .valid_o_gather_pe              (gather_valid_o_4_11),
    .data_o_gather_pe               (gather_data_o_4_11),
    .ready_i_gather_pe              (gather_ready_i_4_11),

    .credit_upd                     (credit_upd[4][11])
);


network_interface #(
    .cast_out                       (cast_out_4_12),
    .gather_out                     (gather_out_4_12),
    .cast_sid                       (cast_sid_4_12),
    .gather_sid                     (gather_sid_4_12)
)ni_4_12(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[4][12]),
    .data_i_cast_nw                 (data_o_cast_nw[4][12]),
    .ready_o_cast_nw                (ready_i_cast_nw[4][12]),
    .valid_o_cast_nw                (valid_i_cast_nw[4][12]),
    .data_o_cast_nw                 (data_i_cast_nw[4][12]),
    .ready_i_cast_nw                (ready_o_cast_nw[4][12]),

    .valid_i_gather_nw              (valid_o_gather_nw[4][12]),
    .data_i_gather_nw               (data_o_gather_nw[4][12]),
    .ready_o_gather_nw              (ready_i_gather_nw[4][12]),
    .valid_o_gather_nw              (valid_i_gather_nw[4][12]),
    .data_o_gather_nw               (data_i_gather_nw[4][12]),
    .ready_i_gather_nw              (ready_o_gather_nw[4][12]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[4][12]),
    .data_i_merge_nw                (data_o_merge_nw[4][12]),
    .ready_o_merge_nw               (ready_i_merge_nw[4][12]),
    .valid_o_merge_nw               (valid_i_merge_nw[4][12]),
    .data_o_merge_nw                (data_i_merge_nw[4][12]),
    .ready_i_merge_nw               (ready_o_merge_nw[4][12]),

    .valid_i_cast_pe                (cast_valid_i_4_12),
    .data_i_cast_pe                 (cast_data_i_4_12),
    .ready_o_cast_pe                (cast_ready_o_4_12),
    .valid_o_cast_pe                (cast_valid_o_4_12),
    .data_o_cast_pe                 (cast_data_o_4_12),
    .ready_i_cast_pe                (cast_ready_i_4_12),

    .valid_i_merge_pe               (merge_valid_i_4_12),
    .data_i_merge_pe                (merge_data_i_4_12),
    .ready_o_merge_pe               (merge_ready_o_4_12),
    .valid_o_merge_pe               (merge_valid_o_4_12),
    .data_o_merge_pe                (merge_data_o_4_12),
    .ready_i_merge_pe               (merge_ready_i_4_12),

    .valid_i_gather_pe              (gather_valid_i_4_12),
    .data_i_gather_pe               (gather_data_i_4_12),
    .ready_o_gather_pe              (gather_ready_o_4_12),
    .valid_o_gather_pe              (gather_valid_o_4_12),
    .data_o_gather_pe               (gather_data_o_4_12),
    .ready_i_gather_pe              (gather_ready_i_4_12),

    .credit_upd                     (credit_upd[4][12])
);


network_interface #(
    .cast_out                       (cast_out_4_13),
    .gather_out                     (gather_out_4_13),
    .cast_sid                       (cast_sid_4_13),
    .gather_sid                     (gather_sid_4_13)
)ni_4_13(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[4][13]),
    .data_i_cast_nw                 (data_o_cast_nw[4][13]),
    .ready_o_cast_nw                (ready_i_cast_nw[4][13]),
    .valid_o_cast_nw                (valid_i_cast_nw[4][13]),
    .data_o_cast_nw                 (data_i_cast_nw[4][13]),
    .ready_i_cast_nw                (ready_o_cast_nw[4][13]),

    .valid_i_gather_nw              (valid_o_gather_nw[4][13]),
    .data_i_gather_nw               (data_o_gather_nw[4][13]),
    .ready_o_gather_nw              (ready_i_gather_nw[4][13]),
    .valid_o_gather_nw              (valid_i_gather_nw[4][13]),
    .data_o_gather_nw               (data_i_gather_nw[4][13]),
    .ready_i_gather_nw              (ready_o_gather_nw[4][13]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[4][13]),
    .data_i_merge_nw                (data_o_merge_nw[4][13]),
    .ready_o_merge_nw               (ready_i_merge_nw[4][13]),
    .valid_o_merge_nw               (valid_i_merge_nw[4][13]),
    .data_o_merge_nw                (data_i_merge_nw[4][13]),
    .ready_i_merge_nw               (ready_o_merge_nw[4][13]),

    .valid_i_cast_pe                (cast_valid_i_4_13),
    .data_i_cast_pe                 (cast_data_i_4_13),
    .ready_o_cast_pe                (cast_ready_o_4_13),
    .valid_o_cast_pe                (cast_valid_o_4_13),
    .data_o_cast_pe                 (cast_data_o_4_13),
    .ready_i_cast_pe                (cast_ready_i_4_13),

    .valid_i_merge_pe               (merge_valid_i_4_13),
    .data_i_merge_pe                (merge_data_i_4_13),
    .ready_o_merge_pe               (merge_ready_o_4_13),
    .valid_o_merge_pe               (merge_valid_o_4_13),
    .data_o_merge_pe                (merge_data_o_4_13),
    .ready_i_merge_pe               (merge_ready_i_4_13),

    .valid_i_gather_pe              (gather_valid_i_4_13),
    .data_i_gather_pe               (gather_data_i_4_13),
    .ready_o_gather_pe              (gather_ready_o_4_13),
    .valid_o_gather_pe              (gather_valid_o_4_13),
    .data_o_gather_pe               (gather_data_o_4_13),
    .ready_i_gather_pe              (gather_ready_i_4_13),

    .credit_upd                     (credit_upd[4][13])
);


network_interface #(
    .cast_out                       (cast_out_4_14),
    .gather_out                     (gather_out_4_14),
    .cast_sid                       (cast_sid_4_14),
    .gather_sid                     (gather_sid_4_14)
)ni_4_14(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[4][14]),
    .data_i_cast_nw                 (data_o_cast_nw[4][14]),
    .ready_o_cast_nw                (ready_i_cast_nw[4][14]),
    .valid_o_cast_nw                (valid_i_cast_nw[4][14]),
    .data_o_cast_nw                 (data_i_cast_nw[4][14]),
    .ready_i_cast_nw                (ready_o_cast_nw[4][14]),

    .valid_i_gather_nw              (valid_o_gather_nw[4][14]),
    .data_i_gather_nw               (data_o_gather_nw[4][14]),
    .ready_o_gather_nw              (ready_i_gather_nw[4][14]),
    .valid_o_gather_nw              (valid_i_gather_nw[4][14]),
    .data_o_gather_nw               (data_i_gather_nw[4][14]),
    .ready_i_gather_nw              (ready_o_gather_nw[4][14]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[4][14]),
    .data_i_merge_nw                (data_o_merge_nw[4][14]),
    .ready_o_merge_nw               (ready_i_merge_nw[4][14]),
    .valid_o_merge_nw               (valid_i_merge_nw[4][14]),
    .data_o_merge_nw                (data_i_merge_nw[4][14]),
    .ready_i_merge_nw               (ready_o_merge_nw[4][14]),

    .valid_i_cast_pe                (cast_valid_i_4_14),
    .data_i_cast_pe                 (cast_data_i_4_14),
    .ready_o_cast_pe                (cast_ready_o_4_14),
    .valid_o_cast_pe                (cast_valid_o_4_14),
    .data_o_cast_pe                 (cast_data_o_4_14),
    .ready_i_cast_pe                (cast_ready_i_4_14),

    .valid_i_merge_pe               (merge_valid_i_4_14),
    .data_i_merge_pe                (merge_data_i_4_14),
    .ready_o_merge_pe               (merge_ready_o_4_14),
    .valid_o_merge_pe               (merge_valid_o_4_14),
    .data_o_merge_pe                (merge_data_o_4_14),
    .ready_i_merge_pe               (merge_ready_i_4_14),

    .valid_i_gather_pe              (gather_valid_i_4_14),
    .data_i_gather_pe               (gather_data_i_4_14),
    .ready_o_gather_pe              (gather_ready_o_4_14),
    .valid_o_gather_pe              (gather_valid_o_4_14),
    .data_o_gather_pe               (gather_data_o_4_14),
    .ready_i_gather_pe              (gather_ready_i_4_14),

    .credit_upd                     (credit_upd[4][14])
);


network_interface #(
    .cast_out                       (cast_out_4_15),
    .gather_out                     (gather_out_4_15),
    .cast_sid                       (cast_sid_4_15),
    .gather_sid                     (gather_sid_4_15)
)ni_4_15(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[4][15]),
    .data_i_cast_nw                 (data_o_cast_nw[4][15]),
    .ready_o_cast_nw                (ready_i_cast_nw[4][15]),
    .valid_o_cast_nw                (valid_i_cast_nw[4][15]),
    .data_o_cast_nw                 (data_i_cast_nw[4][15]),
    .ready_i_cast_nw                (ready_o_cast_nw[4][15]),

    .valid_i_gather_nw              (valid_o_gather_nw[4][15]),
    .data_i_gather_nw               (data_o_gather_nw[4][15]),
    .ready_o_gather_nw              (ready_i_gather_nw[4][15]),
    .valid_o_gather_nw              (valid_i_gather_nw[4][15]),
    .data_o_gather_nw               (data_i_gather_nw[4][15]),
    .ready_i_gather_nw              (ready_o_gather_nw[4][15]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[4][15]),
    .data_i_merge_nw                (data_o_merge_nw[4][15]),
    .ready_o_merge_nw               (ready_i_merge_nw[4][15]),
    .valid_o_merge_nw               (valid_i_merge_nw[4][15]),
    .data_o_merge_nw                (data_i_merge_nw[4][15]),
    .ready_i_merge_nw               (ready_o_merge_nw[4][15]),

    .valid_i_cast_pe                (cast_valid_i_4_15),
    .data_i_cast_pe                 (cast_data_i_4_15),
    .ready_o_cast_pe                (cast_ready_o_4_15),
    .valid_o_cast_pe                (cast_valid_o_4_15),
    .data_o_cast_pe                 (cast_data_o_4_15),
    .ready_i_cast_pe                (cast_ready_i_4_15),

    .valid_i_merge_pe               (merge_valid_i_4_15),
    .data_i_merge_pe                (merge_data_i_4_15),
    .ready_o_merge_pe               (merge_ready_o_4_15),
    .valid_o_merge_pe               (merge_valid_o_4_15),
    .data_o_merge_pe                (merge_data_o_4_15),
    .ready_i_merge_pe               (merge_ready_i_4_15),

    .valid_i_gather_pe              (gather_valid_i_4_15),
    .data_i_gather_pe               (gather_data_i_4_15),
    .ready_o_gather_pe              (gather_ready_o_4_15),
    .valid_o_gather_pe              (gather_valid_o_4_15),
    .data_o_gather_pe               (gather_data_o_4_15),
    .ready_i_gather_pe              (gather_ready_i_4_15),

    .credit_upd                     (credit_upd[4][15])
);


network_interface #(
    .cast_out                       (cast_out_4_16),
    .gather_out                     (gather_out_4_16),
    .cast_sid                       (cast_sid_4_16),
    .gather_sid                     (gather_sid_4_16)
)ni_4_16(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[4][16]),
    .data_i_cast_nw                 (data_o_cast_nw[4][16]),
    .ready_o_cast_nw                (ready_i_cast_nw[4][16]),
    .valid_o_cast_nw                (valid_i_cast_nw[4][16]),
    .data_o_cast_nw                 (data_i_cast_nw[4][16]),
    .ready_i_cast_nw                (ready_o_cast_nw[4][16]),

    .valid_i_gather_nw              (valid_o_gather_nw[4][16]),
    .data_i_gather_nw               (data_o_gather_nw[4][16]),
    .ready_o_gather_nw              (ready_i_gather_nw[4][16]),
    .valid_o_gather_nw              (valid_i_gather_nw[4][16]),
    .data_o_gather_nw               (data_i_gather_nw[4][16]),
    .ready_i_gather_nw              (ready_o_gather_nw[4][16]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[4][16]),
    .data_i_merge_nw                (data_o_merge_nw[4][16]),
    .ready_o_merge_nw               (ready_i_merge_nw[4][16]),
    .valid_o_merge_nw               (valid_i_merge_nw[4][16]),
    .data_o_merge_nw                (data_i_merge_nw[4][16]),
    .ready_i_merge_nw               (ready_o_merge_nw[4][16]),

    .valid_i_cast_pe                (cast_valid_i_4_16),
    .data_i_cast_pe                 (cast_data_i_4_16),
    .ready_o_cast_pe                (cast_ready_o_4_16),
    .valid_o_cast_pe                (cast_valid_o_4_16),
    .data_o_cast_pe                 (cast_data_o_4_16),
    .ready_i_cast_pe                (cast_ready_i_4_16),

    .valid_i_merge_pe               (merge_valid_i_4_16),
    .data_i_merge_pe                (merge_data_i_4_16),
    .ready_o_merge_pe               (merge_ready_o_4_16),
    .valid_o_merge_pe               (merge_valid_o_4_16),
    .data_o_merge_pe                (merge_data_o_4_16),
    .ready_i_merge_pe               (merge_ready_i_4_16),

    .valid_i_gather_pe              (gather_valid_i_4_16),
    .data_i_gather_pe               (gather_data_i_4_16),
    .ready_o_gather_pe              (gather_ready_o_4_16),
    .valid_o_gather_pe              (gather_valid_o_4_16),
    .data_o_gather_pe               (gather_data_o_4_16),
    .ready_i_gather_pe              (gather_ready_i_4_16),

    .credit_upd                     (credit_upd[4][16])
);


network_interface #(
    .cast_out                       (cast_out_4_17),
    .gather_out                     (gather_out_4_17),
    .cast_sid                       (cast_sid_4_17),
    .gather_sid                     (gather_sid_4_17)
)ni_4_17(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[4][17]),
    .data_i_cast_nw                 (data_o_cast_nw[4][17]),
    .ready_o_cast_nw                (ready_i_cast_nw[4][17]),
    .valid_o_cast_nw                (valid_i_cast_nw[4][17]),
    .data_o_cast_nw                 (data_i_cast_nw[4][17]),
    .ready_i_cast_nw                (ready_o_cast_nw[4][17]),

    .valid_i_gather_nw              (valid_o_gather_nw[4][17]),
    .data_i_gather_nw               (data_o_gather_nw[4][17]),
    .ready_o_gather_nw              (ready_i_gather_nw[4][17]),
    .valid_o_gather_nw              (valid_i_gather_nw[4][17]),
    .data_o_gather_nw               (data_i_gather_nw[4][17]),
    .ready_i_gather_nw              (ready_o_gather_nw[4][17]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[4][17]),
    .data_i_merge_nw                (data_o_merge_nw[4][17]),
    .ready_o_merge_nw               (ready_i_merge_nw[4][17]),
    .valid_o_merge_nw               (valid_i_merge_nw[4][17]),
    .data_o_merge_nw                (data_i_merge_nw[4][17]),
    .ready_i_merge_nw               (ready_o_merge_nw[4][17]),

    .valid_i_cast_pe                (cast_valid_i_4_17),
    .data_i_cast_pe                 (cast_data_i_4_17),
    .ready_o_cast_pe                (cast_ready_o_4_17),
    .valid_o_cast_pe                (cast_valid_o_4_17),
    .data_o_cast_pe                 (cast_data_o_4_17),
    .ready_i_cast_pe                (cast_ready_i_4_17),

    .valid_i_merge_pe               (merge_valid_i_4_17),
    .data_i_merge_pe                (merge_data_i_4_17),
    .ready_o_merge_pe               (merge_ready_o_4_17),
    .valid_o_merge_pe               (merge_valid_o_4_17),
    .data_o_merge_pe                (merge_data_o_4_17),
    .ready_i_merge_pe               (merge_ready_i_4_17),

    .valid_i_gather_pe              (gather_valid_i_4_17),
    .data_i_gather_pe               (gather_data_i_4_17),
    .ready_o_gather_pe              (gather_ready_o_4_17),
    .valid_o_gather_pe              (gather_valid_o_4_17),
    .data_o_gather_pe               (gather_data_o_4_17),
    .ready_i_gather_pe              (gather_ready_i_4_17),

    .credit_upd                     (credit_upd[4][17])
);


network_interface #(
    .cast_out                       (cast_out_4_18),
    .gather_out                     (gather_out_4_18),
    .cast_sid                       (cast_sid_4_18),
    .gather_sid                     (gather_sid_4_18)
)ni_4_18(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[4][18]),
    .data_i_cast_nw                 (data_o_cast_nw[4][18]),
    .ready_o_cast_nw                (ready_i_cast_nw[4][18]),
    .valid_o_cast_nw                (valid_i_cast_nw[4][18]),
    .data_o_cast_nw                 (data_i_cast_nw[4][18]),
    .ready_i_cast_nw                (ready_o_cast_nw[4][18]),

    .valid_i_gather_nw              (valid_o_gather_nw[4][18]),
    .data_i_gather_nw               (data_o_gather_nw[4][18]),
    .ready_o_gather_nw              (ready_i_gather_nw[4][18]),
    .valid_o_gather_nw              (valid_i_gather_nw[4][18]),
    .data_o_gather_nw               (data_i_gather_nw[4][18]),
    .ready_i_gather_nw              (ready_o_gather_nw[4][18]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[4][18]),
    .data_i_merge_nw                (data_o_merge_nw[4][18]),
    .ready_o_merge_nw               (ready_i_merge_nw[4][18]),
    .valid_o_merge_nw               (valid_i_merge_nw[4][18]),
    .data_o_merge_nw                (data_i_merge_nw[4][18]),
    .ready_i_merge_nw               (ready_o_merge_nw[4][18]),

    .valid_i_cast_pe                (cast_valid_i_4_18),
    .data_i_cast_pe                 (cast_data_i_4_18),
    .ready_o_cast_pe                (cast_ready_o_4_18),
    .valid_o_cast_pe                (cast_valid_o_4_18),
    .data_o_cast_pe                 (cast_data_o_4_18),
    .ready_i_cast_pe                (cast_ready_i_4_18),

    .valid_i_merge_pe               (merge_valid_i_4_18),
    .data_i_merge_pe                (merge_data_i_4_18),
    .ready_o_merge_pe               (merge_ready_o_4_18),
    .valid_o_merge_pe               (merge_valid_o_4_18),
    .data_o_merge_pe                (merge_data_o_4_18),
    .ready_i_merge_pe               (merge_ready_i_4_18),

    .valid_i_gather_pe              (gather_valid_i_4_18),
    .data_i_gather_pe               (gather_data_i_4_18),
    .ready_o_gather_pe              (gather_ready_o_4_18),
    .valid_o_gather_pe              (gather_valid_o_4_18),
    .data_o_gather_pe               (gather_data_o_4_18),
    .ready_i_gather_pe              (gather_ready_i_4_18),

    .credit_upd                     (credit_upd[4][18])
);


network_interface #(
    .cast_out                       (cast_out_4_19),
    .gather_out                     (gather_out_4_19),
    .cast_sid                       (cast_sid_4_19),
    .gather_sid                     (gather_sid_4_19)
)ni_4_19(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[4][19]),
    .data_i_cast_nw                 (data_o_cast_nw[4][19]),
    .ready_o_cast_nw                (ready_i_cast_nw[4][19]),
    .valid_o_cast_nw                (valid_i_cast_nw[4][19]),
    .data_o_cast_nw                 (data_i_cast_nw[4][19]),
    .ready_i_cast_nw                (ready_o_cast_nw[4][19]),

    .valid_i_gather_nw              (valid_o_gather_nw[4][19]),
    .data_i_gather_nw               (data_o_gather_nw[4][19]),
    .ready_o_gather_nw              (ready_i_gather_nw[4][19]),
    .valid_o_gather_nw              (valid_i_gather_nw[4][19]),
    .data_o_gather_nw               (data_i_gather_nw[4][19]),
    .ready_i_gather_nw              (ready_o_gather_nw[4][19]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[4][19]),
    .data_i_merge_nw                (data_o_merge_nw[4][19]),
    .ready_o_merge_nw               (ready_i_merge_nw[4][19]),
    .valid_o_merge_nw               (valid_i_merge_nw[4][19]),
    .data_o_merge_nw                (data_i_merge_nw[4][19]),
    .ready_i_merge_nw               (ready_o_merge_nw[4][19]),

    .valid_i_cast_pe                (cast_valid_i_4_19),
    .data_i_cast_pe                 (cast_data_i_4_19),
    .ready_o_cast_pe                (cast_ready_o_4_19),
    .valid_o_cast_pe                (cast_valid_o_4_19),
    .data_o_cast_pe                 (cast_data_o_4_19),
    .ready_i_cast_pe                (cast_ready_i_4_19),

    .valid_i_merge_pe               (merge_valid_i_4_19),
    .data_i_merge_pe                (merge_data_i_4_19),
    .ready_o_merge_pe               (merge_ready_o_4_19),
    .valid_o_merge_pe               (merge_valid_o_4_19),
    .data_o_merge_pe                (merge_data_o_4_19),
    .ready_i_merge_pe               (merge_ready_i_4_19),

    .valid_i_gather_pe              (gather_valid_i_4_19),
    .data_i_gather_pe               (gather_data_i_4_19),
    .ready_o_gather_pe              (gather_ready_o_4_19),
    .valid_o_gather_pe              (gather_valid_o_4_19),
    .data_o_gather_pe               (gather_data_o_4_19),
    .ready_i_gather_pe              (gather_ready_i_4_19),

    .credit_upd                     (credit_upd[4][19])
);


network_interface #(
    .cast_out                       (cast_out_4_20),
    .gather_out                     (gather_out_4_20),
    .cast_sid                       (cast_sid_4_20),
    .gather_sid                     (gather_sid_4_20)
)ni_4_20(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[4][20]),
    .data_i_cast_nw                 (data_o_cast_nw[4][20]),
    .ready_o_cast_nw                (ready_i_cast_nw[4][20]),
    .valid_o_cast_nw                (valid_i_cast_nw[4][20]),
    .data_o_cast_nw                 (data_i_cast_nw[4][20]),
    .ready_i_cast_nw                (ready_o_cast_nw[4][20]),

    .valid_i_gather_nw              (valid_o_gather_nw[4][20]),
    .data_i_gather_nw               (data_o_gather_nw[4][20]),
    .ready_o_gather_nw              (ready_i_gather_nw[4][20]),
    .valid_o_gather_nw              (valid_i_gather_nw[4][20]),
    .data_o_gather_nw               (data_i_gather_nw[4][20]),
    .ready_i_gather_nw              (ready_o_gather_nw[4][20]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[4][20]),
    .data_i_merge_nw                (data_o_merge_nw[4][20]),
    .ready_o_merge_nw               (ready_i_merge_nw[4][20]),
    .valid_o_merge_nw               (valid_i_merge_nw[4][20]),
    .data_o_merge_nw                (data_i_merge_nw[4][20]),
    .ready_i_merge_nw               (ready_o_merge_nw[4][20]),

    .valid_i_cast_pe                (cast_valid_i_4_20),
    .data_i_cast_pe                 (cast_data_i_4_20),
    .ready_o_cast_pe                (cast_ready_o_4_20),
    .valid_o_cast_pe                (cast_valid_o_4_20),
    .data_o_cast_pe                 (cast_data_o_4_20),
    .ready_i_cast_pe                (cast_ready_i_4_20),

    .valid_i_merge_pe               (merge_valid_i_4_20),
    .data_i_merge_pe                (merge_data_i_4_20),
    .ready_o_merge_pe               (merge_ready_o_4_20),
    .valid_o_merge_pe               (merge_valid_o_4_20),
    .data_o_merge_pe                (merge_data_o_4_20),
    .ready_i_merge_pe               (merge_ready_i_4_20),

    .valid_i_gather_pe              (gather_valid_i_4_20),
    .data_i_gather_pe               (gather_data_i_4_20),
    .ready_o_gather_pe              (gather_ready_o_4_20),
    .valid_o_gather_pe              (gather_valid_o_4_20),
    .data_o_gather_pe               (gather_data_o_4_20),
    .ready_i_gather_pe              (gather_ready_i_4_20),

    .credit_upd                     (credit_upd[4][20])
);


network_interface #(
    .cast_out                       (cast_out_4_21),
    .gather_out                     (gather_out_4_21),
    .cast_sid                       (cast_sid_4_21),
    .gather_sid                     (gather_sid_4_21)
)ni_4_21(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[4][21]),
    .data_i_cast_nw                 (data_o_cast_nw[4][21]),
    .ready_o_cast_nw                (ready_i_cast_nw[4][21]),
    .valid_o_cast_nw                (valid_i_cast_nw[4][21]),
    .data_o_cast_nw                 (data_i_cast_nw[4][21]),
    .ready_i_cast_nw                (ready_o_cast_nw[4][21]),

    .valid_i_gather_nw              (valid_o_gather_nw[4][21]),
    .data_i_gather_nw               (data_o_gather_nw[4][21]),
    .ready_o_gather_nw              (ready_i_gather_nw[4][21]),
    .valid_o_gather_nw              (valid_i_gather_nw[4][21]),
    .data_o_gather_nw               (data_i_gather_nw[4][21]),
    .ready_i_gather_nw              (ready_o_gather_nw[4][21]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[4][21]),
    .data_i_merge_nw                (data_o_merge_nw[4][21]),
    .ready_o_merge_nw               (ready_i_merge_nw[4][21]),
    .valid_o_merge_nw               (valid_i_merge_nw[4][21]),
    .data_o_merge_nw                (data_i_merge_nw[4][21]),
    .ready_i_merge_nw               (ready_o_merge_nw[4][21]),

    .valid_i_cast_pe                (cast_valid_i_4_21),
    .data_i_cast_pe                 (cast_data_i_4_21),
    .ready_o_cast_pe                (cast_ready_o_4_21),
    .valid_o_cast_pe                (cast_valid_o_4_21),
    .data_o_cast_pe                 (cast_data_o_4_21),
    .ready_i_cast_pe                (cast_ready_i_4_21),

    .valid_i_merge_pe               (merge_valid_i_4_21),
    .data_i_merge_pe                (merge_data_i_4_21),
    .ready_o_merge_pe               (merge_ready_o_4_21),
    .valid_o_merge_pe               (merge_valid_o_4_21),
    .data_o_merge_pe                (merge_data_o_4_21),
    .ready_i_merge_pe               (merge_ready_i_4_21),

    .valid_i_gather_pe              (gather_valid_i_4_21),
    .data_i_gather_pe               (gather_data_i_4_21),
    .ready_o_gather_pe              (gather_ready_o_4_21),
    .valid_o_gather_pe              (gather_valid_o_4_21),
    .data_o_gather_pe               (gather_data_o_4_21),
    .ready_i_gather_pe              (gather_ready_i_4_21),

    .credit_upd                     (credit_upd[4][21])
);


network_interface #(
    .cast_out                       (cast_out_4_22),
    .gather_out                     (gather_out_4_22),
    .cast_sid                       (cast_sid_4_22),
    .gather_sid                     (gather_sid_4_22)
)ni_4_22(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[4][22]),
    .data_i_cast_nw                 (data_o_cast_nw[4][22]),
    .ready_o_cast_nw                (ready_i_cast_nw[4][22]),
    .valid_o_cast_nw                (valid_i_cast_nw[4][22]),
    .data_o_cast_nw                 (data_i_cast_nw[4][22]),
    .ready_i_cast_nw                (ready_o_cast_nw[4][22]),

    .valid_i_gather_nw              (valid_o_gather_nw[4][22]),
    .data_i_gather_nw               (data_o_gather_nw[4][22]),
    .ready_o_gather_nw              (ready_i_gather_nw[4][22]),
    .valid_o_gather_nw              (valid_i_gather_nw[4][22]),
    .data_o_gather_nw               (data_i_gather_nw[4][22]),
    .ready_i_gather_nw              (ready_o_gather_nw[4][22]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[4][22]),
    .data_i_merge_nw                (data_o_merge_nw[4][22]),
    .ready_o_merge_nw               (ready_i_merge_nw[4][22]),
    .valid_o_merge_nw               (valid_i_merge_nw[4][22]),
    .data_o_merge_nw                (data_i_merge_nw[4][22]),
    .ready_i_merge_nw               (ready_o_merge_nw[4][22]),

    .valid_i_cast_pe                (cast_valid_i_4_22),
    .data_i_cast_pe                 (cast_data_i_4_22),
    .ready_o_cast_pe                (cast_ready_o_4_22),
    .valid_o_cast_pe                (cast_valid_o_4_22),
    .data_o_cast_pe                 (cast_data_o_4_22),
    .ready_i_cast_pe                (cast_ready_i_4_22),

    .valid_i_merge_pe               (merge_valid_i_4_22),
    .data_i_merge_pe                (merge_data_i_4_22),
    .ready_o_merge_pe               (merge_ready_o_4_22),
    .valid_o_merge_pe               (merge_valid_o_4_22),
    .data_o_merge_pe                (merge_data_o_4_22),
    .ready_i_merge_pe               (merge_ready_i_4_22),

    .valid_i_gather_pe              (gather_valid_i_4_22),
    .data_i_gather_pe               (gather_data_i_4_22),
    .ready_o_gather_pe              (gather_ready_o_4_22),
    .valid_o_gather_pe              (gather_valid_o_4_22),
    .data_o_gather_pe               (gather_data_o_4_22),
    .ready_i_gather_pe              (gather_ready_i_4_22),

    .credit_upd                     (credit_upd[4][22])
);


network_interface #(
    .cast_out                       (cast_out_4_23),
    .gather_out                     (gather_out_4_23),
    .cast_sid                       (cast_sid_4_23),
    .gather_sid                     (gather_sid_4_23)
)ni_4_23(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[4][23]),
    .data_i_cast_nw                 (data_o_cast_nw[4][23]),
    .ready_o_cast_nw                (ready_i_cast_nw[4][23]),
    .valid_o_cast_nw                (valid_i_cast_nw[4][23]),
    .data_o_cast_nw                 (data_i_cast_nw[4][23]),
    .ready_i_cast_nw                (ready_o_cast_nw[4][23]),

    .valid_i_gather_nw              (valid_o_gather_nw[4][23]),
    .data_i_gather_nw               (data_o_gather_nw[4][23]),
    .ready_o_gather_nw              (ready_i_gather_nw[4][23]),
    .valid_o_gather_nw              (valid_i_gather_nw[4][23]),
    .data_o_gather_nw               (data_i_gather_nw[4][23]),
    .ready_i_gather_nw              (ready_o_gather_nw[4][23]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[4][23]),
    .data_i_merge_nw                (data_o_merge_nw[4][23]),
    .ready_o_merge_nw               (ready_i_merge_nw[4][23]),
    .valid_o_merge_nw               (valid_i_merge_nw[4][23]),
    .data_o_merge_nw                (data_i_merge_nw[4][23]),
    .ready_i_merge_nw               (ready_o_merge_nw[4][23]),

    .valid_i_cast_pe                (cast_valid_i_4_23),
    .data_i_cast_pe                 (cast_data_i_4_23),
    .ready_o_cast_pe                (cast_ready_o_4_23),
    .valid_o_cast_pe                (cast_valid_o_4_23),
    .data_o_cast_pe                 (cast_data_o_4_23),
    .ready_i_cast_pe                (cast_ready_i_4_23),

    .valid_i_merge_pe               (merge_valid_i_4_23),
    .data_i_merge_pe                (merge_data_i_4_23),
    .ready_o_merge_pe               (merge_ready_o_4_23),
    .valid_o_merge_pe               (merge_valid_o_4_23),
    .data_o_merge_pe                (merge_data_o_4_23),
    .ready_i_merge_pe               (merge_ready_i_4_23),

    .valid_i_gather_pe              (gather_valid_i_4_23),
    .data_i_gather_pe               (gather_data_i_4_23),
    .ready_o_gather_pe              (gather_ready_o_4_23),
    .valid_o_gather_pe              (gather_valid_o_4_23),
    .data_o_gather_pe               (gather_data_o_4_23),
    .ready_i_gather_pe              (gather_ready_i_4_23),

    .credit_upd                     (credit_upd[4][23])
);


network_interface #(
    .cast_out                       (cast_out_4_24),
    .gather_out                     (gather_out_4_24),
    .cast_sid                       (cast_sid_4_24),
    .gather_sid                     (gather_sid_4_24)
)ni_4_24(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[4][24]),
    .data_i_cast_nw                 (data_o_cast_nw[4][24]),
    .ready_o_cast_nw                (ready_i_cast_nw[4][24]),
    .valid_o_cast_nw                (valid_i_cast_nw[4][24]),
    .data_o_cast_nw                 (data_i_cast_nw[4][24]),
    .ready_i_cast_nw                (ready_o_cast_nw[4][24]),

    .valid_i_gather_nw              (valid_o_gather_nw[4][24]),
    .data_i_gather_nw               (data_o_gather_nw[4][24]),
    .ready_o_gather_nw              (ready_i_gather_nw[4][24]),
    .valid_o_gather_nw              (valid_i_gather_nw[4][24]),
    .data_o_gather_nw               (data_i_gather_nw[4][24]),
    .ready_i_gather_nw              (ready_o_gather_nw[4][24]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[4][24]),
    .data_i_merge_nw                (data_o_merge_nw[4][24]),
    .ready_o_merge_nw               (ready_i_merge_nw[4][24]),
    .valid_o_merge_nw               (valid_i_merge_nw[4][24]),
    .data_o_merge_nw                (data_i_merge_nw[4][24]),
    .ready_i_merge_nw               (ready_o_merge_nw[4][24]),

    .valid_i_cast_pe                (cast_valid_i_4_24),
    .data_i_cast_pe                 (cast_data_i_4_24),
    .ready_o_cast_pe                (cast_ready_o_4_24),
    .valid_o_cast_pe                (cast_valid_o_4_24),
    .data_o_cast_pe                 (cast_data_o_4_24),
    .ready_i_cast_pe                (cast_ready_i_4_24),

    .valid_i_merge_pe               (merge_valid_i_4_24),
    .data_i_merge_pe                (merge_data_i_4_24),
    .ready_o_merge_pe               (merge_ready_o_4_24),
    .valid_o_merge_pe               (merge_valid_o_4_24),
    .data_o_merge_pe                (merge_data_o_4_24),
    .ready_i_merge_pe               (merge_ready_i_4_24),

    .valid_i_gather_pe              (gather_valid_i_4_24),
    .data_i_gather_pe               (gather_data_i_4_24),
    .ready_o_gather_pe              (gather_ready_o_4_24),
    .valid_o_gather_pe              (gather_valid_o_4_24),
    .data_o_gather_pe               (gather_data_o_4_24),
    .ready_i_gather_pe              (gather_ready_i_4_24),

    .credit_upd                     (credit_upd[4][24])
);


network_interface #(
    .cast_out                       (cast_out_5_0),
    .gather_out                     (gather_out_5_0),
    .cast_sid                       (cast_sid_5_0),
    .gather_sid                     (gather_sid_5_0)
)ni_5_0(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[5][0]),
    .data_i_cast_nw                 (data_o_cast_nw[5][0]),
    .ready_o_cast_nw                (ready_i_cast_nw[5][0]),
    .valid_o_cast_nw                (valid_i_cast_nw[5][0]),
    .data_o_cast_nw                 (data_i_cast_nw[5][0]),
    .ready_i_cast_nw                (ready_o_cast_nw[5][0]),

    .valid_i_gather_nw              (valid_o_gather_nw[5][0]),
    .data_i_gather_nw               (data_o_gather_nw[5][0]),
    .ready_o_gather_nw              (ready_i_gather_nw[5][0]),
    .valid_o_gather_nw              (valid_i_gather_nw[5][0]),
    .data_o_gather_nw               (data_i_gather_nw[5][0]),
    .ready_i_gather_nw              (ready_o_gather_nw[5][0]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[5][0]),
    .data_i_merge_nw                (data_o_merge_nw[5][0]),
    .ready_o_merge_nw               (ready_i_merge_nw[5][0]),
    .valid_o_merge_nw               (valid_i_merge_nw[5][0]),
    .data_o_merge_nw                (data_i_merge_nw[5][0]),
    .ready_i_merge_nw               (ready_o_merge_nw[5][0]),

    .valid_i_cast_pe                (cast_valid_i_5_0),
    .data_i_cast_pe                 (cast_data_i_5_0),
    .ready_o_cast_pe                (cast_ready_o_5_0),
    .valid_o_cast_pe                (cast_valid_o_5_0),
    .data_o_cast_pe                 (cast_data_o_5_0),
    .ready_i_cast_pe                (cast_ready_i_5_0),

    .valid_i_merge_pe               (merge_valid_i_5_0),
    .data_i_merge_pe                (merge_data_i_5_0),
    .ready_o_merge_pe               (merge_ready_o_5_0),
    .valid_o_merge_pe               (merge_valid_o_5_0),
    .data_o_merge_pe                (merge_data_o_5_0),
    .ready_i_merge_pe               (merge_ready_i_5_0),

    .valid_i_gather_pe              (gather_valid_i_5_0),
    .data_i_gather_pe               (gather_data_i_5_0),
    .ready_o_gather_pe              (gather_ready_o_5_0),
    .valid_o_gather_pe              (gather_valid_o_5_0),
    .data_o_gather_pe               (gather_data_o_5_0),
    .ready_i_gather_pe              (gather_ready_i_5_0),

    .credit_upd                     (credit_upd[5][0])
);


network_interface #(
    .cast_out                       (cast_out_5_1),
    .gather_out                     (gather_out_5_1),
    .cast_sid                       (cast_sid_5_1),
    .gather_sid                     (gather_sid_5_1)
)ni_5_1(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[5][1]),
    .data_i_cast_nw                 (data_o_cast_nw[5][1]),
    .ready_o_cast_nw                (ready_i_cast_nw[5][1]),
    .valid_o_cast_nw                (valid_i_cast_nw[5][1]),
    .data_o_cast_nw                 (data_i_cast_nw[5][1]),
    .ready_i_cast_nw                (ready_o_cast_nw[5][1]),

    .valid_i_gather_nw              (valid_o_gather_nw[5][1]),
    .data_i_gather_nw               (data_o_gather_nw[5][1]),
    .ready_o_gather_nw              (ready_i_gather_nw[5][1]),
    .valid_o_gather_nw              (valid_i_gather_nw[5][1]),
    .data_o_gather_nw               (data_i_gather_nw[5][1]),
    .ready_i_gather_nw              (ready_o_gather_nw[5][1]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[5][1]),
    .data_i_merge_nw                (data_o_merge_nw[5][1]),
    .ready_o_merge_nw               (ready_i_merge_nw[5][1]),
    .valid_o_merge_nw               (valid_i_merge_nw[5][1]),
    .data_o_merge_nw                (data_i_merge_nw[5][1]),
    .ready_i_merge_nw               (ready_o_merge_nw[5][1]),

    .valid_i_cast_pe                (cast_valid_i_5_1),
    .data_i_cast_pe                 (cast_data_i_5_1),
    .ready_o_cast_pe                (cast_ready_o_5_1),
    .valid_o_cast_pe                (cast_valid_o_5_1),
    .data_o_cast_pe                 (cast_data_o_5_1),
    .ready_i_cast_pe                (cast_ready_i_5_1),

    .valid_i_merge_pe               (merge_valid_i_5_1),
    .data_i_merge_pe                (merge_data_i_5_1),
    .ready_o_merge_pe               (merge_ready_o_5_1),
    .valid_o_merge_pe               (merge_valid_o_5_1),
    .data_o_merge_pe                (merge_data_o_5_1),
    .ready_i_merge_pe               (merge_ready_i_5_1),

    .valid_i_gather_pe              (gather_valid_i_5_1),
    .data_i_gather_pe               (gather_data_i_5_1),
    .ready_o_gather_pe              (gather_ready_o_5_1),
    .valid_o_gather_pe              (gather_valid_o_5_1),
    .data_o_gather_pe               (gather_data_o_5_1),
    .ready_i_gather_pe              (gather_ready_i_5_1),

    .credit_upd                     (credit_upd[5][1])
);


network_interface #(
    .cast_out                       (cast_out_5_2),
    .gather_out                     (gather_out_5_2),
    .cast_sid                       (cast_sid_5_2),
    .gather_sid                     (gather_sid_5_2)
)ni_5_2(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[5][2]),
    .data_i_cast_nw                 (data_o_cast_nw[5][2]),
    .ready_o_cast_nw                (ready_i_cast_nw[5][2]),
    .valid_o_cast_nw                (valid_i_cast_nw[5][2]),
    .data_o_cast_nw                 (data_i_cast_nw[5][2]),
    .ready_i_cast_nw                (ready_o_cast_nw[5][2]),

    .valid_i_gather_nw              (valid_o_gather_nw[5][2]),
    .data_i_gather_nw               (data_o_gather_nw[5][2]),
    .ready_o_gather_nw              (ready_i_gather_nw[5][2]),
    .valid_o_gather_nw              (valid_i_gather_nw[5][2]),
    .data_o_gather_nw               (data_i_gather_nw[5][2]),
    .ready_i_gather_nw              (ready_o_gather_nw[5][2]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[5][2]),
    .data_i_merge_nw                (data_o_merge_nw[5][2]),
    .ready_o_merge_nw               (ready_i_merge_nw[5][2]),
    .valid_o_merge_nw               (valid_i_merge_nw[5][2]),
    .data_o_merge_nw                (data_i_merge_nw[5][2]),
    .ready_i_merge_nw               (ready_o_merge_nw[5][2]),

    .valid_i_cast_pe                (cast_valid_i_5_2),
    .data_i_cast_pe                 (cast_data_i_5_2),
    .ready_o_cast_pe                (cast_ready_o_5_2),
    .valid_o_cast_pe                (cast_valid_o_5_2),
    .data_o_cast_pe                 (cast_data_o_5_2),
    .ready_i_cast_pe                (cast_ready_i_5_2),

    .valid_i_merge_pe               (merge_valid_i_5_2),
    .data_i_merge_pe                (merge_data_i_5_2),
    .ready_o_merge_pe               (merge_ready_o_5_2),
    .valid_o_merge_pe               (merge_valid_o_5_2),
    .data_o_merge_pe                (merge_data_o_5_2),
    .ready_i_merge_pe               (merge_ready_i_5_2),

    .valid_i_gather_pe              (gather_valid_i_5_2),
    .data_i_gather_pe               (gather_data_i_5_2),
    .ready_o_gather_pe              (gather_ready_o_5_2),
    .valid_o_gather_pe              (gather_valid_o_5_2),
    .data_o_gather_pe               (gather_data_o_5_2),
    .ready_i_gather_pe              (gather_ready_i_5_2),

    .credit_upd                     (credit_upd[5][2])
);


network_interface #(
    .cast_out                       (cast_out_5_3),
    .gather_out                     (gather_out_5_3),
    .cast_sid                       (cast_sid_5_3),
    .gather_sid                     (gather_sid_5_3)
)ni_5_3(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[5][3]),
    .data_i_cast_nw                 (data_o_cast_nw[5][3]),
    .ready_o_cast_nw                (ready_i_cast_nw[5][3]),
    .valid_o_cast_nw                (valid_i_cast_nw[5][3]),
    .data_o_cast_nw                 (data_i_cast_nw[5][3]),
    .ready_i_cast_nw                (ready_o_cast_nw[5][3]),

    .valid_i_gather_nw              (valid_o_gather_nw[5][3]),
    .data_i_gather_nw               (data_o_gather_nw[5][3]),
    .ready_o_gather_nw              (ready_i_gather_nw[5][3]),
    .valid_o_gather_nw              (valid_i_gather_nw[5][3]),
    .data_o_gather_nw               (data_i_gather_nw[5][3]),
    .ready_i_gather_nw              (ready_o_gather_nw[5][3]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[5][3]),
    .data_i_merge_nw                (data_o_merge_nw[5][3]),
    .ready_o_merge_nw               (ready_i_merge_nw[5][3]),
    .valid_o_merge_nw               (valid_i_merge_nw[5][3]),
    .data_o_merge_nw                (data_i_merge_nw[5][3]),
    .ready_i_merge_nw               (ready_o_merge_nw[5][3]),

    .valid_i_cast_pe                (cast_valid_i_5_3),
    .data_i_cast_pe                 (cast_data_i_5_3),
    .ready_o_cast_pe                (cast_ready_o_5_3),
    .valid_o_cast_pe                (cast_valid_o_5_3),
    .data_o_cast_pe                 (cast_data_o_5_3),
    .ready_i_cast_pe                (cast_ready_i_5_3),

    .valid_i_merge_pe               (merge_valid_i_5_3),
    .data_i_merge_pe                (merge_data_i_5_3),
    .ready_o_merge_pe               (merge_ready_o_5_3),
    .valid_o_merge_pe               (merge_valid_o_5_3),
    .data_o_merge_pe                (merge_data_o_5_3),
    .ready_i_merge_pe               (merge_ready_i_5_3),

    .valid_i_gather_pe              (gather_valid_i_5_3),
    .data_i_gather_pe               (gather_data_i_5_3),
    .ready_o_gather_pe              (gather_ready_o_5_3),
    .valid_o_gather_pe              (gather_valid_o_5_3),
    .data_o_gather_pe               (gather_data_o_5_3),
    .ready_i_gather_pe              (gather_ready_i_5_3),

    .credit_upd                     (credit_upd[5][3])
);


network_interface #(
    .cast_out                       (cast_out_5_4),
    .gather_out                     (gather_out_5_4),
    .cast_sid                       (cast_sid_5_4),
    .gather_sid                     (gather_sid_5_4)
)ni_5_4(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[5][4]),
    .data_i_cast_nw                 (data_o_cast_nw[5][4]),
    .ready_o_cast_nw                (ready_i_cast_nw[5][4]),
    .valid_o_cast_nw                (valid_i_cast_nw[5][4]),
    .data_o_cast_nw                 (data_i_cast_nw[5][4]),
    .ready_i_cast_nw                (ready_o_cast_nw[5][4]),

    .valid_i_gather_nw              (valid_o_gather_nw[5][4]),
    .data_i_gather_nw               (data_o_gather_nw[5][4]),
    .ready_o_gather_nw              (ready_i_gather_nw[5][4]),
    .valid_o_gather_nw              (valid_i_gather_nw[5][4]),
    .data_o_gather_nw               (data_i_gather_nw[5][4]),
    .ready_i_gather_nw              (ready_o_gather_nw[5][4]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[5][4]),
    .data_i_merge_nw                (data_o_merge_nw[5][4]),
    .ready_o_merge_nw               (ready_i_merge_nw[5][4]),
    .valid_o_merge_nw               (valid_i_merge_nw[5][4]),
    .data_o_merge_nw                (data_i_merge_nw[5][4]),
    .ready_i_merge_nw               (ready_o_merge_nw[5][4]),

    .valid_i_cast_pe                (cast_valid_i_5_4),
    .data_i_cast_pe                 (cast_data_i_5_4),
    .ready_o_cast_pe                (cast_ready_o_5_4),
    .valid_o_cast_pe                (cast_valid_o_5_4),
    .data_o_cast_pe                 (cast_data_o_5_4),
    .ready_i_cast_pe                (cast_ready_i_5_4),

    .valid_i_merge_pe               (merge_valid_i_5_4),
    .data_i_merge_pe                (merge_data_i_5_4),
    .ready_o_merge_pe               (merge_ready_o_5_4),
    .valid_o_merge_pe               (merge_valid_o_5_4),
    .data_o_merge_pe                (merge_data_o_5_4),
    .ready_i_merge_pe               (merge_ready_i_5_4),

    .valid_i_gather_pe              (gather_valid_i_5_4),
    .data_i_gather_pe               (gather_data_i_5_4),
    .ready_o_gather_pe              (gather_ready_o_5_4),
    .valid_o_gather_pe              (gather_valid_o_5_4),
    .data_o_gather_pe               (gather_data_o_5_4),
    .ready_i_gather_pe              (gather_ready_i_5_4),

    .credit_upd                     (credit_upd[5][4])
);


network_interface #(
    .cast_out                       (cast_out_5_5),
    .gather_out                     (gather_out_5_5),
    .cast_sid                       (cast_sid_5_5),
    .gather_sid                     (gather_sid_5_5)
)ni_5_5(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[5][5]),
    .data_i_cast_nw                 (data_o_cast_nw[5][5]),
    .ready_o_cast_nw                (ready_i_cast_nw[5][5]),
    .valid_o_cast_nw                (valid_i_cast_nw[5][5]),
    .data_o_cast_nw                 (data_i_cast_nw[5][5]),
    .ready_i_cast_nw                (ready_o_cast_nw[5][5]),

    .valid_i_gather_nw              (valid_o_gather_nw[5][5]),
    .data_i_gather_nw               (data_o_gather_nw[5][5]),
    .ready_o_gather_nw              (ready_i_gather_nw[5][5]),
    .valid_o_gather_nw              (valid_i_gather_nw[5][5]),
    .data_o_gather_nw               (data_i_gather_nw[5][5]),
    .ready_i_gather_nw              (ready_o_gather_nw[5][5]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[5][5]),
    .data_i_merge_nw                (data_o_merge_nw[5][5]),
    .ready_o_merge_nw               (ready_i_merge_nw[5][5]),
    .valid_o_merge_nw               (valid_i_merge_nw[5][5]),
    .data_o_merge_nw                (data_i_merge_nw[5][5]),
    .ready_i_merge_nw               (ready_o_merge_nw[5][5]),

    .valid_i_cast_pe                (cast_valid_i_5_5),
    .data_i_cast_pe                 (cast_data_i_5_5),
    .ready_o_cast_pe                (cast_ready_o_5_5),
    .valid_o_cast_pe                (cast_valid_o_5_5),
    .data_o_cast_pe                 (cast_data_o_5_5),
    .ready_i_cast_pe                (cast_ready_i_5_5),

    .valid_i_merge_pe               (merge_valid_i_5_5),
    .data_i_merge_pe                (merge_data_i_5_5),
    .ready_o_merge_pe               (merge_ready_o_5_5),
    .valid_o_merge_pe               (merge_valid_o_5_5),
    .data_o_merge_pe                (merge_data_o_5_5),
    .ready_i_merge_pe               (merge_ready_i_5_5),

    .valid_i_gather_pe              (gather_valid_i_5_5),
    .data_i_gather_pe               (gather_data_i_5_5),
    .ready_o_gather_pe              (gather_ready_o_5_5),
    .valid_o_gather_pe              (gather_valid_o_5_5),
    .data_o_gather_pe               (gather_data_o_5_5),
    .ready_i_gather_pe              (gather_ready_i_5_5),

    .credit_upd                     (credit_upd[5][5])
);


network_interface #(
    .cast_out                       (cast_out_5_6),
    .gather_out                     (gather_out_5_6),
    .cast_sid                       (cast_sid_5_6),
    .gather_sid                     (gather_sid_5_6)
)ni_5_6(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[5][6]),
    .data_i_cast_nw                 (data_o_cast_nw[5][6]),
    .ready_o_cast_nw                (ready_i_cast_nw[5][6]),
    .valid_o_cast_nw                (valid_i_cast_nw[5][6]),
    .data_o_cast_nw                 (data_i_cast_nw[5][6]),
    .ready_i_cast_nw                (ready_o_cast_nw[5][6]),

    .valid_i_gather_nw              (valid_o_gather_nw[5][6]),
    .data_i_gather_nw               (data_o_gather_nw[5][6]),
    .ready_o_gather_nw              (ready_i_gather_nw[5][6]),
    .valid_o_gather_nw              (valid_i_gather_nw[5][6]),
    .data_o_gather_nw               (data_i_gather_nw[5][6]),
    .ready_i_gather_nw              (ready_o_gather_nw[5][6]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[5][6]),
    .data_i_merge_nw                (data_o_merge_nw[5][6]),
    .ready_o_merge_nw               (ready_i_merge_nw[5][6]),
    .valid_o_merge_nw               (valid_i_merge_nw[5][6]),
    .data_o_merge_nw                (data_i_merge_nw[5][6]),
    .ready_i_merge_nw               (ready_o_merge_nw[5][6]),

    .valid_i_cast_pe                (cast_valid_i_5_6),
    .data_i_cast_pe                 (cast_data_i_5_6),
    .ready_o_cast_pe                (cast_ready_o_5_6),
    .valid_o_cast_pe                (cast_valid_o_5_6),
    .data_o_cast_pe                 (cast_data_o_5_6),
    .ready_i_cast_pe                (cast_ready_i_5_6),

    .valid_i_merge_pe               (merge_valid_i_5_6),
    .data_i_merge_pe                (merge_data_i_5_6),
    .ready_o_merge_pe               (merge_ready_o_5_6),
    .valid_o_merge_pe               (merge_valid_o_5_6),
    .data_o_merge_pe                (merge_data_o_5_6),
    .ready_i_merge_pe               (merge_ready_i_5_6),

    .valid_i_gather_pe              (gather_valid_i_5_6),
    .data_i_gather_pe               (gather_data_i_5_6),
    .ready_o_gather_pe              (gather_ready_o_5_6),
    .valid_o_gather_pe              (gather_valid_o_5_6),
    .data_o_gather_pe               (gather_data_o_5_6),
    .ready_i_gather_pe              (gather_ready_i_5_6),

    .credit_upd                     (credit_upd[5][6])
);


network_interface #(
    .cast_out                       (cast_out_5_7),
    .gather_out                     (gather_out_5_7),
    .cast_sid                       (cast_sid_5_7),
    .gather_sid                     (gather_sid_5_7)
)ni_5_7(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[5][7]),
    .data_i_cast_nw                 (data_o_cast_nw[5][7]),
    .ready_o_cast_nw                (ready_i_cast_nw[5][7]),
    .valid_o_cast_nw                (valid_i_cast_nw[5][7]),
    .data_o_cast_nw                 (data_i_cast_nw[5][7]),
    .ready_i_cast_nw                (ready_o_cast_nw[5][7]),

    .valid_i_gather_nw              (valid_o_gather_nw[5][7]),
    .data_i_gather_nw               (data_o_gather_nw[5][7]),
    .ready_o_gather_nw              (ready_i_gather_nw[5][7]),
    .valid_o_gather_nw              (valid_i_gather_nw[5][7]),
    .data_o_gather_nw               (data_i_gather_nw[5][7]),
    .ready_i_gather_nw              (ready_o_gather_nw[5][7]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[5][7]),
    .data_i_merge_nw                (data_o_merge_nw[5][7]),
    .ready_o_merge_nw               (ready_i_merge_nw[5][7]),
    .valid_o_merge_nw               (valid_i_merge_nw[5][7]),
    .data_o_merge_nw                (data_i_merge_nw[5][7]),
    .ready_i_merge_nw               (ready_o_merge_nw[5][7]),

    .valid_i_cast_pe                (cast_valid_i_5_7),
    .data_i_cast_pe                 (cast_data_i_5_7),
    .ready_o_cast_pe                (cast_ready_o_5_7),
    .valid_o_cast_pe                (cast_valid_o_5_7),
    .data_o_cast_pe                 (cast_data_o_5_7),
    .ready_i_cast_pe                (cast_ready_i_5_7),

    .valid_i_merge_pe               (merge_valid_i_5_7),
    .data_i_merge_pe                (merge_data_i_5_7),
    .ready_o_merge_pe               (merge_ready_o_5_7),
    .valid_o_merge_pe               (merge_valid_o_5_7),
    .data_o_merge_pe                (merge_data_o_5_7),
    .ready_i_merge_pe               (merge_ready_i_5_7),

    .valid_i_gather_pe              (gather_valid_i_5_7),
    .data_i_gather_pe               (gather_data_i_5_7),
    .ready_o_gather_pe              (gather_ready_o_5_7),
    .valid_o_gather_pe              (gather_valid_o_5_7),
    .data_o_gather_pe               (gather_data_o_5_7),
    .ready_i_gather_pe              (gather_ready_i_5_7),

    .credit_upd                     (credit_upd[5][7])
);


network_interface #(
    .cast_out                       (cast_out_5_8),
    .gather_out                     (gather_out_5_8),
    .cast_sid                       (cast_sid_5_8),
    .gather_sid                     (gather_sid_5_8)
)ni_5_8(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[5][8]),
    .data_i_cast_nw                 (data_o_cast_nw[5][8]),
    .ready_o_cast_nw                (ready_i_cast_nw[5][8]),
    .valid_o_cast_nw                (valid_i_cast_nw[5][8]),
    .data_o_cast_nw                 (data_i_cast_nw[5][8]),
    .ready_i_cast_nw                (ready_o_cast_nw[5][8]),

    .valid_i_gather_nw              (valid_o_gather_nw[5][8]),
    .data_i_gather_nw               (data_o_gather_nw[5][8]),
    .ready_o_gather_nw              (ready_i_gather_nw[5][8]),
    .valid_o_gather_nw              (valid_i_gather_nw[5][8]),
    .data_o_gather_nw               (data_i_gather_nw[5][8]),
    .ready_i_gather_nw              (ready_o_gather_nw[5][8]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[5][8]),
    .data_i_merge_nw                (data_o_merge_nw[5][8]),
    .ready_o_merge_nw               (ready_i_merge_nw[5][8]),
    .valid_o_merge_nw               (valid_i_merge_nw[5][8]),
    .data_o_merge_nw                (data_i_merge_nw[5][8]),
    .ready_i_merge_nw               (ready_o_merge_nw[5][8]),

    .valid_i_cast_pe                (cast_valid_i_5_8),
    .data_i_cast_pe                 (cast_data_i_5_8),
    .ready_o_cast_pe                (cast_ready_o_5_8),
    .valid_o_cast_pe                (cast_valid_o_5_8),
    .data_o_cast_pe                 (cast_data_o_5_8),
    .ready_i_cast_pe                (cast_ready_i_5_8),

    .valid_i_merge_pe               (merge_valid_i_5_8),
    .data_i_merge_pe                (merge_data_i_5_8),
    .ready_o_merge_pe               (merge_ready_o_5_8),
    .valid_o_merge_pe               (merge_valid_o_5_8),
    .data_o_merge_pe                (merge_data_o_5_8),
    .ready_i_merge_pe               (merge_ready_i_5_8),

    .valid_i_gather_pe              (gather_valid_i_5_8),
    .data_i_gather_pe               (gather_data_i_5_8),
    .ready_o_gather_pe              (gather_ready_o_5_8),
    .valid_o_gather_pe              (gather_valid_o_5_8),
    .data_o_gather_pe               (gather_data_o_5_8),
    .ready_i_gather_pe              (gather_ready_i_5_8),

    .credit_upd                     (credit_upd[5][8])
);


network_interface #(
    .cast_out                       (cast_out_5_9),
    .gather_out                     (gather_out_5_9),
    .cast_sid                       (cast_sid_5_9),
    .gather_sid                     (gather_sid_5_9)
)ni_5_9(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[5][9]),
    .data_i_cast_nw                 (data_o_cast_nw[5][9]),
    .ready_o_cast_nw                (ready_i_cast_nw[5][9]),
    .valid_o_cast_nw                (valid_i_cast_nw[5][9]),
    .data_o_cast_nw                 (data_i_cast_nw[5][9]),
    .ready_i_cast_nw                (ready_o_cast_nw[5][9]),

    .valid_i_gather_nw              (valid_o_gather_nw[5][9]),
    .data_i_gather_nw               (data_o_gather_nw[5][9]),
    .ready_o_gather_nw              (ready_i_gather_nw[5][9]),
    .valid_o_gather_nw              (valid_i_gather_nw[5][9]),
    .data_o_gather_nw               (data_i_gather_nw[5][9]),
    .ready_i_gather_nw              (ready_o_gather_nw[5][9]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[5][9]),
    .data_i_merge_nw                (data_o_merge_nw[5][9]),
    .ready_o_merge_nw               (ready_i_merge_nw[5][9]),
    .valid_o_merge_nw               (valid_i_merge_nw[5][9]),
    .data_o_merge_nw                (data_i_merge_nw[5][9]),
    .ready_i_merge_nw               (ready_o_merge_nw[5][9]),

    .valid_i_cast_pe                (cast_valid_i_5_9),
    .data_i_cast_pe                 (cast_data_i_5_9),
    .ready_o_cast_pe                (cast_ready_o_5_9),
    .valid_o_cast_pe                (cast_valid_o_5_9),
    .data_o_cast_pe                 (cast_data_o_5_9),
    .ready_i_cast_pe                (cast_ready_i_5_9),

    .valid_i_merge_pe               (merge_valid_i_5_9),
    .data_i_merge_pe                (merge_data_i_5_9),
    .ready_o_merge_pe               (merge_ready_o_5_9),
    .valid_o_merge_pe               (merge_valid_o_5_9),
    .data_o_merge_pe                (merge_data_o_5_9),
    .ready_i_merge_pe               (merge_ready_i_5_9),

    .valid_i_gather_pe              (gather_valid_i_5_9),
    .data_i_gather_pe               (gather_data_i_5_9),
    .ready_o_gather_pe              (gather_ready_o_5_9),
    .valid_o_gather_pe              (gather_valid_o_5_9),
    .data_o_gather_pe               (gather_data_o_5_9),
    .ready_i_gather_pe              (gather_ready_i_5_9),

    .credit_upd                     (credit_upd[5][9])
);


network_interface #(
    .cast_out                       (cast_out_5_10),
    .gather_out                     (gather_out_5_10),
    .cast_sid                       (cast_sid_5_10),
    .gather_sid                     (gather_sid_5_10)
)ni_5_10(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[5][10]),
    .data_i_cast_nw                 (data_o_cast_nw[5][10]),
    .ready_o_cast_nw                (ready_i_cast_nw[5][10]),
    .valid_o_cast_nw                (valid_i_cast_nw[5][10]),
    .data_o_cast_nw                 (data_i_cast_nw[5][10]),
    .ready_i_cast_nw                (ready_o_cast_nw[5][10]),

    .valid_i_gather_nw              (valid_o_gather_nw[5][10]),
    .data_i_gather_nw               (data_o_gather_nw[5][10]),
    .ready_o_gather_nw              (ready_i_gather_nw[5][10]),
    .valid_o_gather_nw              (valid_i_gather_nw[5][10]),
    .data_o_gather_nw               (data_i_gather_nw[5][10]),
    .ready_i_gather_nw              (ready_o_gather_nw[5][10]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[5][10]),
    .data_i_merge_nw                (data_o_merge_nw[5][10]),
    .ready_o_merge_nw               (ready_i_merge_nw[5][10]),
    .valid_o_merge_nw               (valid_i_merge_nw[5][10]),
    .data_o_merge_nw                (data_i_merge_nw[5][10]),
    .ready_i_merge_nw               (ready_o_merge_nw[5][10]),

    .valid_i_cast_pe                (cast_valid_i_5_10),
    .data_i_cast_pe                 (cast_data_i_5_10),
    .ready_o_cast_pe                (cast_ready_o_5_10),
    .valid_o_cast_pe                (cast_valid_o_5_10),
    .data_o_cast_pe                 (cast_data_o_5_10),
    .ready_i_cast_pe                (cast_ready_i_5_10),

    .valid_i_merge_pe               (merge_valid_i_5_10),
    .data_i_merge_pe                (merge_data_i_5_10),
    .ready_o_merge_pe               (merge_ready_o_5_10),
    .valid_o_merge_pe               (merge_valid_o_5_10),
    .data_o_merge_pe                (merge_data_o_5_10),
    .ready_i_merge_pe               (merge_ready_i_5_10),

    .valid_i_gather_pe              (gather_valid_i_5_10),
    .data_i_gather_pe               (gather_data_i_5_10),
    .ready_o_gather_pe              (gather_ready_o_5_10),
    .valid_o_gather_pe              (gather_valid_o_5_10),
    .data_o_gather_pe               (gather_data_o_5_10),
    .ready_i_gather_pe              (gather_ready_i_5_10),

    .credit_upd                     (credit_upd[5][10])
);


network_interface #(
    .cast_out                       (cast_out_5_11),
    .gather_out                     (gather_out_5_11),
    .cast_sid                       (cast_sid_5_11),
    .gather_sid                     (gather_sid_5_11)
)ni_5_11(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[5][11]),
    .data_i_cast_nw                 (data_o_cast_nw[5][11]),
    .ready_o_cast_nw                (ready_i_cast_nw[5][11]),
    .valid_o_cast_nw                (valid_i_cast_nw[5][11]),
    .data_o_cast_nw                 (data_i_cast_nw[5][11]),
    .ready_i_cast_nw                (ready_o_cast_nw[5][11]),

    .valid_i_gather_nw              (valid_o_gather_nw[5][11]),
    .data_i_gather_nw               (data_o_gather_nw[5][11]),
    .ready_o_gather_nw              (ready_i_gather_nw[5][11]),
    .valid_o_gather_nw              (valid_i_gather_nw[5][11]),
    .data_o_gather_nw               (data_i_gather_nw[5][11]),
    .ready_i_gather_nw              (ready_o_gather_nw[5][11]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[5][11]),
    .data_i_merge_nw                (data_o_merge_nw[5][11]),
    .ready_o_merge_nw               (ready_i_merge_nw[5][11]),
    .valid_o_merge_nw               (valid_i_merge_nw[5][11]),
    .data_o_merge_nw                (data_i_merge_nw[5][11]),
    .ready_i_merge_nw               (ready_o_merge_nw[5][11]),

    .valid_i_cast_pe                (cast_valid_i_5_11),
    .data_i_cast_pe                 (cast_data_i_5_11),
    .ready_o_cast_pe                (cast_ready_o_5_11),
    .valid_o_cast_pe                (cast_valid_o_5_11),
    .data_o_cast_pe                 (cast_data_o_5_11),
    .ready_i_cast_pe                (cast_ready_i_5_11),

    .valid_i_merge_pe               (merge_valid_i_5_11),
    .data_i_merge_pe                (merge_data_i_5_11),
    .ready_o_merge_pe               (merge_ready_o_5_11),
    .valid_o_merge_pe               (merge_valid_o_5_11),
    .data_o_merge_pe                (merge_data_o_5_11),
    .ready_i_merge_pe               (merge_ready_i_5_11),

    .valid_i_gather_pe              (gather_valid_i_5_11),
    .data_i_gather_pe               (gather_data_i_5_11),
    .ready_o_gather_pe              (gather_ready_o_5_11),
    .valid_o_gather_pe              (gather_valid_o_5_11),
    .data_o_gather_pe               (gather_data_o_5_11),
    .ready_i_gather_pe              (gather_ready_i_5_11),

    .credit_upd                     (credit_upd[5][11])
);


network_interface #(
    .cast_out                       (cast_out_5_12),
    .gather_out                     (gather_out_5_12),
    .cast_sid                       (cast_sid_5_12),
    .gather_sid                     (gather_sid_5_12)
)ni_5_12(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[5][12]),
    .data_i_cast_nw                 (data_o_cast_nw[5][12]),
    .ready_o_cast_nw                (ready_i_cast_nw[5][12]),
    .valid_o_cast_nw                (valid_i_cast_nw[5][12]),
    .data_o_cast_nw                 (data_i_cast_nw[5][12]),
    .ready_i_cast_nw                (ready_o_cast_nw[5][12]),

    .valid_i_gather_nw              (valid_o_gather_nw[5][12]),
    .data_i_gather_nw               (data_o_gather_nw[5][12]),
    .ready_o_gather_nw              (ready_i_gather_nw[5][12]),
    .valid_o_gather_nw              (valid_i_gather_nw[5][12]),
    .data_o_gather_nw               (data_i_gather_nw[5][12]),
    .ready_i_gather_nw              (ready_o_gather_nw[5][12]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[5][12]),
    .data_i_merge_nw                (data_o_merge_nw[5][12]),
    .ready_o_merge_nw               (ready_i_merge_nw[5][12]),
    .valid_o_merge_nw               (valid_i_merge_nw[5][12]),
    .data_o_merge_nw                (data_i_merge_nw[5][12]),
    .ready_i_merge_nw               (ready_o_merge_nw[5][12]),

    .valid_i_cast_pe                (cast_valid_i_5_12),
    .data_i_cast_pe                 (cast_data_i_5_12),
    .ready_o_cast_pe                (cast_ready_o_5_12),
    .valid_o_cast_pe                (cast_valid_o_5_12),
    .data_o_cast_pe                 (cast_data_o_5_12),
    .ready_i_cast_pe                (cast_ready_i_5_12),

    .valid_i_merge_pe               (merge_valid_i_5_12),
    .data_i_merge_pe                (merge_data_i_5_12),
    .ready_o_merge_pe               (merge_ready_o_5_12),
    .valid_o_merge_pe               (merge_valid_o_5_12),
    .data_o_merge_pe                (merge_data_o_5_12),
    .ready_i_merge_pe               (merge_ready_i_5_12),

    .valid_i_gather_pe              (gather_valid_i_5_12),
    .data_i_gather_pe               (gather_data_i_5_12),
    .ready_o_gather_pe              (gather_ready_o_5_12),
    .valid_o_gather_pe              (gather_valid_o_5_12),
    .data_o_gather_pe               (gather_data_o_5_12),
    .ready_i_gather_pe              (gather_ready_i_5_12),

    .credit_upd                     (credit_upd[5][12])
);


network_interface #(
    .cast_out                       (cast_out_5_13),
    .gather_out                     (gather_out_5_13),
    .cast_sid                       (cast_sid_5_13),
    .gather_sid                     (gather_sid_5_13)
)ni_5_13(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[5][13]),
    .data_i_cast_nw                 (data_o_cast_nw[5][13]),
    .ready_o_cast_nw                (ready_i_cast_nw[5][13]),
    .valid_o_cast_nw                (valid_i_cast_nw[5][13]),
    .data_o_cast_nw                 (data_i_cast_nw[5][13]),
    .ready_i_cast_nw                (ready_o_cast_nw[5][13]),

    .valid_i_gather_nw              (valid_o_gather_nw[5][13]),
    .data_i_gather_nw               (data_o_gather_nw[5][13]),
    .ready_o_gather_nw              (ready_i_gather_nw[5][13]),
    .valid_o_gather_nw              (valid_i_gather_nw[5][13]),
    .data_o_gather_nw               (data_i_gather_nw[5][13]),
    .ready_i_gather_nw              (ready_o_gather_nw[5][13]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[5][13]),
    .data_i_merge_nw                (data_o_merge_nw[5][13]),
    .ready_o_merge_nw               (ready_i_merge_nw[5][13]),
    .valid_o_merge_nw               (valid_i_merge_nw[5][13]),
    .data_o_merge_nw                (data_i_merge_nw[5][13]),
    .ready_i_merge_nw               (ready_o_merge_nw[5][13]),

    .valid_i_cast_pe                (cast_valid_i_5_13),
    .data_i_cast_pe                 (cast_data_i_5_13),
    .ready_o_cast_pe                (cast_ready_o_5_13),
    .valid_o_cast_pe                (cast_valid_o_5_13),
    .data_o_cast_pe                 (cast_data_o_5_13),
    .ready_i_cast_pe                (cast_ready_i_5_13),

    .valid_i_merge_pe               (merge_valid_i_5_13),
    .data_i_merge_pe                (merge_data_i_5_13),
    .ready_o_merge_pe               (merge_ready_o_5_13),
    .valid_o_merge_pe               (merge_valid_o_5_13),
    .data_o_merge_pe                (merge_data_o_5_13),
    .ready_i_merge_pe               (merge_ready_i_5_13),

    .valid_i_gather_pe              (gather_valid_i_5_13),
    .data_i_gather_pe               (gather_data_i_5_13),
    .ready_o_gather_pe              (gather_ready_o_5_13),
    .valid_o_gather_pe              (gather_valid_o_5_13),
    .data_o_gather_pe               (gather_data_o_5_13),
    .ready_i_gather_pe              (gather_ready_i_5_13),

    .credit_upd                     (credit_upd[5][13])
);


network_interface #(
    .cast_out                       (cast_out_5_14),
    .gather_out                     (gather_out_5_14),
    .cast_sid                       (cast_sid_5_14),
    .gather_sid                     (gather_sid_5_14)
)ni_5_14(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[5][14]),
    .data_i_cast_nw                 (data_o_cast_nw[5][14]),
    .ready_o_cast_nw                (ready_i_cast_nw[5][14]),
    .valid_o_cast_nw                (valid_i_cast_nw[5][14]),
    .data_o_cast_nw                 (data_i_cast_nw[5][14]),
    .ready_i_cast_nw                (ready_o_cast_nw[5][14]),

    .valid_i_gather_nw              (valid_o_gather_nw[5][14]),
    .data_i_gather_nw               (data_o_gather_nw[5][14]),
    .ready_o_gather_nw              (ready_i_gather_nw[5][14]),
    .valid_o_gather_nw              (valid_i_gather_nw[5][14]),
    .data_o_gather_nw               (data_i_gather_nw[5][14]),
    .ready_i_gather_nw              (ready_o_gather_nw[5][14]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[5][14]),
    .data_i_merge_nw                (data_o_merge_nw[5][14]),
    .ready_o_merge_nw               (ready_i_merge_nw[5][14]),
    .valid_o_merge_nw               (valid_i_merge_nw[5][14]),
    .data_o_merge_nw                (data_i_merge_nw[5][14]),
    .ready_i_merge_nw               (ready_o_merge_nw[5][14]),

    .valid_i_cast_pe                (cast_valid_i_5_14),
    .data_i_cast_pe                 (cast_data_i_5_14),
    .ready_o_cast_pe                (cast_ready_o_5_14),
    .valid_o_cast_pe                (cast_valid_o_5_14),
    .data_o_cast_pe                 (cast_data_o_5_14),
    .ready_i_cast_pe                (cast_ready_i_5_14),

    .valid_i_merge_pe               (merge_valid_i_5_14),
    .data_i_merge_pe                (merge_data_i_5_14),
    .ready_o_merge_pe               (merge_ready_o_5_14),
    .valid_o_merge_pe               (merge_valid_o_5_14),
    .data_o_merge_pe                (merge_data_o_5_14),
    .ready_i_merge_pe               (merge_ready_i_5_14),

    .valid_i_gather_pe              (gather_valid_i_5_14),
    .data_i_gather_pe               (gather_data_i_5_14),
    .ready_o_gather_pe              (gather_ready_o_5_14),
    .valid_o_gather_pe              (gather_valid_o_5_14),
    .data_o_gather_pe               (gather_data_o_5_14),
    .ready_i_gather_pe              (gather_ready_i_5_14),

    .credit_upd                     (credit_upd[5][14])
);


network_interface #(
    .cast_out                       (cast_out_5_15),
    .gather_out                     (gather_out_5_15),
    .cast_sid                       (cast_sid_5_15),
    .gather_sid                     (gather_sid_5_15)
)ni_5_15(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[5][15]),
    .data_i_cast_nw                 (data_o_cast_nw[5][15]),
    .ready_o_cast_nw                (ready_i_cast_nw[5][15]),
    .valid_o_cast_nw                (valid_i_cast_nw[5][15]),
    .data_o_cast_nw                 (data_i_cast_nw[5][15]),
    .ready_i_cast_nw                (ready_o_cast_nw[5][15]),

    .valid_i_gather_nw              (valid_o_gather_nw[5][15]),
    .data_i_gather_nw               (data_o_gather_nw[5][15]),
    .ready_o_gather_nw              (ready_i_gather_nw[5][15]),
    .valid_o_gather_nw              (valid_i_gather_nw[5][15]),
    .data_o_gather_nw               (data_i_gather_nw[5][15]),
    .ready_i_gather_nw              (ready_o_gather_nw[5][15]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[5][15]),
    .data_i_merge_nw                (data_o_merge_nw[5][15]),
    .ready_o_merge_nw               (ready_i_merge_nw[5][15]),
    .valid_o_merge_nw               (valid_i_merge_nw[5][15]),
    .data_o_merge_nw                (data_i_merge_nw[5][15]),
    .ready_i_merge_nw               (ready_o_merge_nw[5][15]),

    .valid_i_cast_pe                (cast_valid_i_5_15),
    .data_i_cast_pe                 (cast_data_i_5_15),
    .ready_o_cast_pe                (cast_ready_o_5_15),
    .valid_o_cast_pe                (cast_valid_o_5_15),
    .data_o_cast_pe                 (cast_data_o_5_15),
    .ready_i_cast_pe                (cast_ready_i_5_15),

    .valid_i_merge_pe               (merge_valid_i_5_15),
    .data_i_merge_pe                (merge_data_i_5_15),
    .ready_o_merge_pe               (merge_ready_o_5_15),
    .valid_o_merge_pe               (merge_valid_o_5_15),
    .data_o_merge_pe                (merge_data_o_5_15),
    .ready_i_merge_pe               (merge_ready_i_5_15),

    .valid_i_gather_pe              (gather_valid_i_5_15),
    .data_i_gather_pe               (gather_data_i_5_15),
    .ready_o_gather_pe              (gather_ready_o_5_15),
    .valid_o_gather_pe              (gather_valid_o_5_15),
    .data_o_gather_pe               (gather_data_o_5_15),
    .ready_i_gather_pe              (gather_ready_i_5_15),

    .credit_upd                     (credit_upd[5][15])
);


network_interface #(
    .cast_out                       (cast_out_5_16),
    .gather_out                     (gather_out_5_16),
    .cast_sid                       (cast_sid_5_16),
    .gather_sid                     (gather_sid_5_16)
)ni_5_16(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[5][16]),
    .data_i_cast_nw                 (data_o_cast_nw[5][16]),
    .ready_o_cast_nw                (ready_i_cast_nw[5][16]),
    .valid_o_cast_nw                (valid_i_cast_nw[5][16]),
    .data_o_cast_nw                 (data_i_cast_nw[5][16]),
    .ready_i_cast_nw                (ready_o_cast_nw[5][16]),

    .valid_i_gather_nw              (valid_o_gather_nw[5][16]),
    .data_i_gather_nw               (data_o_gather_nw[5][16]),
    .ready_o_gather_nw              (ready_i_gather_nw[5][16]),
    .valid_o_gather_nw              (valid_i_gather_nw[5][16]),
    .data_o_gather_nw               (data_i_gather_nw[5][16]),
    .ready_i_gather_nw              (ready_o_gather_nw[5][16]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[5][16]),
    .data_i_merge_nw                (data_o_merge_nw[5][16]),
    .ready_o_merge_nw               (ready_i_merge_nw[5][16]),
    .valid_o_merge_nw               (valid_i_merge_nw[5][16]),
    .data_o_merge_nw                (data_i_merge_nw[5][16]),
    .ready_i_merge_nw               (ready_o_merge_nw[5][16]),

    .valid_i_cast_pe                (cast_valid_i_5_16),
    .data_i_cast_pe                 (cast_data_i_5_16),
    .ready_o_cast_pe                (cast_ready_o_5_16),
    .valid_o_cast_pe                (cast_valid_o_5_16),
    .data_o_cast_pe                 (cast_data_o_5_16),
    .ready_i_cast_pe                (cast_ready_i_5_16),

    .valid_i_merge_pe               (merge_valid_i_5_16),
    .data_i_merge_pe                (merge_data_i_5_16),
    .ready_o_merge_pe               (merge_ready_o_5_16),
    .valid_o_merge_pe               (merge_valid_o_5_16),
    .data_o_merge_pe                (merge_data_o_5_16),
    .ready_i_merge_pe               (merge_ready_i_5_16),

    .valid_i_gather_pe              (gather_valid_i_5_16),
    .data_i_gather_pe               (gather_data_i_5_16),
    .ready_o_gather_pe              (gather_ready_o_5_16),
    .valid_o_gather_pe              (gather_valid_o_5_16),
    .data_o_gather_pe               (gather_data_o_5_16),
    .ready_i_gather_pe              (gather_ready_i_5_16),

    .credit_upd                     (credit_upd[5][16])
);


network_interface #(
    .cast_out                       (cast_out_5_17),
    .gather_out                     (gather_out_5_17),
    .cast_sid                       (cast_sid_5_17),
    .gather_sid                     (gather_sid_5_17)
)ni_5_17(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[5][17]),
    .data_i_cast_nw                 (data_o_cast_nw[5][17]),
    .ready_o_cast_nw                (ready_i_cast_nw[5][17]),
    .valid_o_cast_nw                (valid_i_cast_nw[5][17]),
    .data_o_cast_nw                 (data_i_cast_nw[5][17]),
    .ready_i_cast_nw                (ready_o_cast_nw[5][17]),

    .valid_i_gather_nw              (valid_o_gather_nw[5][17]),
    .data_i_gather_nw               (data_o_gather_nw[5][17]),
    .ready_o_gather_nw              (ready_i_gather_nw[5][17]),
    .valid_o_gather_nw              (valid_i_gather_nw[5][17]),
    .data_o_gather_nw               (data_i_gather_nw[5][17]),
    .ready_i_gather_nw              (ready_o_gather_nw[5][17]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[5][17]),
    .data_i_merge_nw                (data_o_merge_nw[5][17]),
    .ready_o_merge_nw               (ready_i_merge_nw[5][17]),
    .valid_o_merge_nw               (valid_i_merge_nw[5][17]),
    .data_o_merge_nw                (data_i_merge_nw[5][17]),
    .ready_i_merge_nw               (ready_o_merge_nw[5][17]),

    .valid_i_cast_pe                (cast_valid_i_5_17),
    .data_i_cast_pe                 (cast_data_i_5_17),
    .ready_o_cast_pe                (cast_ready_o_5_17),
    .valid_o_cast_pe                (cast_valid_o_5_17),
    .data_o_cast_pe                 (cast_data_o_5_17),
    .ready_i_cast_pe                (cast_ready_i_5_17),

    .valid_i_merge_pe               (merge_valid_i_5_17),
    .data_i_merge_pe                (merge_data_i_5_17),
    .ready_o_merge_pe               (merge_ready_o_5_17),
    .valid_o_merge_pe               (merge_valid_o_5_17),
    .data_o_merge_pe                (merge_data_o_5_17),
    .ready_i_merge_pe               (merge_ready_i_5_17),

    .valid_i_gather_pe              (gather_valid_i_5_17),
    .data_i_gather_pe               (gather_data_i_5_17),
    .ready_o_gather_pe              (gather_ready_o_5_17),
    .valid_o_gather_pe              (gather_valid_o_5_17),
    .data_o_gather_pe               (gather_data_o_5_17),
    .ready_i_gather_pe              (gather_ready_i_5_17),

    .credit_upd                     (credit_upd[5][17])
);


network_interface #(
    .cast_out                       (cast_out_5_18),
    .gather_out                     (gather_out_5_18),
    .cast_sid                       (cast_sid_5_18),
    .gather_sid                     (gather_sid_5_18)
)ni_5_18(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[5][18]),
    .data_i_cast_nw                 (data_o_cast_nw[5][18]),
    .ready_o_cast_nw                (ready_i_cast_nw[5][18]),
    .valid_o_cast_nw                (valid_i_cast_nw[5][18]),
    .data_o_cast_nw                 (data_i_cast_nw[5][18]),
    .ready_i_cast_nw                (ready_o_cast_nw[5][18]),

    .valid_i_gather_nw              (valid_o_gather_nw[5][18]),
    .data_i_gather_nw               (data_o_gather_nw[5][18]),
    .ready_o_gather_nw              (ready_i_gather_nw[5][18]),
    .valid_o_gather_nw              (valid_i_gather_nw[5][18]),
    .data_o_gather_nw               (data_i_gather_nw[5][18]),
    .ready_i_gather_nw              (ready_o_gather_nw[5][18]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[5][18]),
    .data_i_merge_nw                (data_o_merge_nw[5][18]),
    .ready_o_merge_nw               (ready_i_merge_nw[5][18]),
    .valid_o_merge_nw               (valid_i_merge_nw[5][18]),
    .data_o_merge_nw                (data_i_merge_nw[5][18]),
    .ready_i_merge_nw               (ready_o_merge_nw[5][18]),

    .valid_i_cast_pe                (cast_valid_i_5_18),
    .data_i_cast_pe                 (cast_data_i_5_18),
    .ready_o_cast_pe                (cast_ready_o_5_18),
    .valid_o_cast_pe                (cast_valid_o_5_18),
    .data_o_cast_pe                 (cast_data_o_5_18),
    .ready_i_cast_pe                (cast_ready_i_5_18),

    .valid_i_merge_pe               (merge_valid_i_5_18),
    .data_i_merge_pe                (merge_data_i_5_18),
    .ready_o_merge_pe               (merge_ready_o_5_18),
    .valid_o_merge_pe               (merge_valid_o_5_18),
    .data_o_merge_pe                (merge_data_o_5_18),
    .ready_i_merge_pe               (merge_ready_i_5_18),

    .valid_i_gather_pe              (gather_valid_i_5_18),
    .data_i_gather_pe               (gather_data_i_5_18),
    .ready_o_gather_pe              (gather_ready_o_5_18),
    .valid_o_gather_pe              (gather_valid_o_5_18),
    .data_o_gather_pe               (gather_data_o_5_18),
    .ready_i_gather_pe              (gather_ready_i_5_18),

    .credit_upd                     (credit_upd[5][18])
);


network_interface #(
    .cast_out                       (cast_out_5_19),
    .gather_out                     (gather_out_5_19),
    .cast_sid                       (cast_sid_5_19),
    .gather_sid                     (gather_sid_5_19)
)ni_5_19(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[5][19]),
    .data_i_cast_nw                 (data_o_cast_nw[5][19]),
    .ready_o_cast_nw                (ready_i_cast_nw[5][19]),
    .valid_o_cast_nw                (valid_i_cast_nw[5][19]),
    .data_o_cast_nw                 (data_i_cast_nw[5][19]),
    .ready_i_cast_nw                (ready_o_cast_nw[5][19]),

    .valid_i_gather_nw              (valid_o_gather_nw[5][19]),
    .data_i_gather_nw               (data_o_gather_nw[5][19]),
    .ready_o_gather_nw              (ready_i_gather_nw[5][19]),
    .valid_o_gather_nw              (valid_i_gather_nw[5][19]),
    .data_o_gather_nw               (data_i_gather_nw[5][19]),
    .ready_i_gather_nw              (ready_o_gather_nw[5][19]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[5][19]),
    .data_i_merge_nw                (data_o_merge_nw[5][19]),
    .ready_o_merge_nw               (ready_i_merge_nw[5][19]),
    .valid_o_merge_nw               (valid_i_merge_nw[5][19]),
    .data_o_merge_nw                (data_i_merge_nw[5][19]),
    .ready_i_merge_nw               (ready_o_merge_nw[5][19]),

    .valid_i_cast_pe                (cast_valid_i_5_19),
    .data_i_cast_pe                 (cast_data_i_5_19),
    .ready_o_cast_pe                (cast_ready_o_5_19),
    .valid_o_cast_pe                (cast_valid_o_5_19),
    .data_o_cast_pe                 (cast_data_o_5_19),
    .ready_i_cast_pe                (cast_ready_i_5_19),

    .valid_i_merge_pe               (merge_valid_i_5_19),
    .data_i_merge_pe                (merge_data_i_5_19),
    .ready_o_merge_pe               (merge_ready_o_5_19),
    .valid_o_merge_pe               (merge_valid_o_5_19),
    .data_o_merge_pe                (merge_data_o_5_19),
    .ready_i_merge_pe               (merge_ready_i_5_19),

    .valid_i_gather_pe              (gather_valid_i_5_19),
    .data_i_gather_pe               (gather_data_i_5_19),
    .ready_o_gather_pe              (gather_ready_o_5_19),
    .valid_o_gather_pe              (gather_valid_o_5_19),
    .data_o_gather_pe               (gather_data_o_5_19),
    .ready_i_gather_pe              (gather_ready_i_5_19),

    .credit_upd                     (credit_upd[5][19])
);


network_interface #(
    .cast_out                       (cast_out_5_20),
    .gather_out                     (gather_out_5_20),
    .cast_sid                       (cast_sid_5_20),
    .gather_sid                     (gather_sid_5_20)
)ni_5_20(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[5][20]),
    .data_i_cast_nw                 (data_o_cast_nw[5][20]),
    .ready_o_cast_nw                (ready_i_cast_nw[5][20]),
    .valid_o_cast_nw                (valid_i_cast_nw[5][20]),
    .data_o_cast_nw                 (data_i_cast_nw[5][20]),
    .ready_i_cast_nw                (ready_o_cast_nw[5][20]),

    .valid_i_gather_nw              (valid_o_gather_nw[5][20]),
    .data_i_gather_nw               (data_o_gather_nw[5][20]),
    .ready_o_gather_nw              (ready_i_gather_nw[5][20]),
    .valid_o_gather_nw              (valid_i_gather_nw[5][20]),
    .data_o_gather_nw               (data_i_gather_nw[5][20]),
    .ready_i_gather_nw              (ready_o_gather_nw[5][20]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[5][20]),
    .data_i_merge_nw                (data_o_merge_nw[5][20]),
    .ready_o_merge_nw               (ready_i_merge_nw[5][20]),
    .valid_o_merge_nw               (valid_i_merge_nw[5][20]),
    .data_o_merge_nw                (data_i_merge_nw[5][20]),
    .ready_i_merge_nw               (ready_o_merge_nw[5][20]),

    .valid_i_cast_pe                (cast_valid_i_5_20),
    .data_i_cast_pe                 (cast_data_i_5_20),
    .ready_o_cast_pe                (cast_ready_o_5_20),
    .valid_o_cast_pe                (cast_valid_o_5_20),
    .data_o_cast_pe                 (cast_data_o_5_20),
    .ready_i_cast_pe                (cast_ready_i_5_20),

    .valid_i_merge_pe               (merge_valid_i_5_20),
    .data_i_merge_pe                (merge_data_i_5_20),
    .ready_o_merge_pe               (merge_ready_o_5_20),
    .valid_o_merge_pe               (merge_valid_o_5_20),
    .data_o_merge_pe                (merge_data_o_5_20),
    .ready_i_merge_pe               (merge_ready_i_5_20),

    .valid_i_gather_pe              (gather_valid_i_5_20),
    .data_i_gather_pe               (gather_data_i_5_20),
    .ready_o_gather_pe              (gather_ready_o_5_20),
    .valid_o_gather_pe              (gather_valid_o_5_20),
    .data_o_gather_pe               (gather_data_o_5_20),
    .ready_i_gather_pe              (gather_ready_i_5_20),

    .credit_upd                     (credit_upd[5][20])
);


network_interface #(
    .cast_out                       (cast_out_5_21),
    .gather_out                     (gather_out_5_21),
    .cast_sid                       (cast_sid_5_21),
    .gather_sid                     (gather_sid_5_21)
)ni_5_21(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[5][21]),
    .data_i_cast_nw                 (data_o_cast_nw[5][21]),
    .ready_o_cast_nw                (ready_i_cast_nw[5][21]),
    .valid_o_cast_nw                (valid_i_cast_nw[5][21]),
    .data_o_cast_nw                 (data_i_cast_nw[5][21]),
    .ready_i_cast_nw                (ready_o_cast_nw[5][21]),

    .valid_i_gather_nw              (valid_o_gather_nw[5][21]),
    .data_i_gather_nw               (data_o_gather_nw[5][21]),
    .ready_o_gather_nw              (ready_i_gather_nw[5][21]),
    .valid_o_gather_nw              (valid_i_gather_nw[5][21]),
    .data_o_gather_nw               (data_i_gather_nw[5][21]),
    .ready_i_gather_nw              (ready_o_gather_nw[5][21]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[5][21]),
    .data_i_merge_nw                (data_o_merge_nw[5][21]),
    .ready_o_merge_nw               (ready_i_merge_nw[5][21]),
    .valid_o_merge_nw               (valid_i_merge_nw[5][21]),
    .data_o_merge_nw                (data_i_merge_nw[5][21]),
    .ready_i_merge_nw               (ready_o_merge_nw[5][21]),

    .valid_i_cast_pe                (cast_valid_i_5_21),
    .data_i_cast_pe                 (cast_data_i_5_21),
    .ready_o_cast_pe                (cast_ready_o_5_21),
    .valid_o_cast_pe                (cast_valid_o_5_21),
    .data_o_cast_pe                 (cast_data_o_5_21),
    .ready_i_cast_pe                (cast_ready_i_5_21),

    .valid_i_merge_pe               (merge_valid_i_5_21),
    .data_i_merge_pe                (merge_data_i_5_21),
    .ready_o_merge_pe               (merge_ready_o_5_21),
    .valid_o_merge_pe               (merge_valid_o_5_21),
    .data_o_merge_pe                (merge_data_o_5_21),
    .ready_i_merge_pe               (merge_ready_i_5_21),

    .valid_i_gather_pe              (gather_valid_i_5_21),
    .data_i_gather_pe               (gather_data_i_5_21),
    .ready_o_gather_pe              (gather_ready_o_5_21),
    .valid_o_gather_pe              (gather_valid_o_5_21),
    .data_o_gather_pe               (gather_data_o_5_21),
    .ready_i_gather_pe              (gather_ready_i_5_21),

    .credit_upd                     (credit_upd[5][21])
);


network_interface #(
    .cast_out                       (cast_out_5_22),
    .gather_out                     (gather_out_5_22),
    .cast_sid                       (cast_sid_5_22),
    .gather_sid                     (gather_sid_5_22)
)ni_5_22(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[5][22]),
    .data_i_cast_nw                 (data_o_cast_nw[5][22]),
    .ready_o_cast_nw                (ready_i_cast_nw[5][22]),
    .valid_o_cast_nw                (valid_i_cast_nw[5][22]),
    .data_o_cast_nw                 (data_i_cast_nw[5][22]),
    .ready_i_cast_nw                (ready_o_cast_nw[5][22]),

    .valid_i_gather_nw              (valid_o_gather_nw[5][22]),
    .data_i_gather_nw               (data_o_gather_nw[5][22]),
    .ready_o_gather_nw              (ready_i_gather_nw[5][22]),
    .valid_o_gather_nw              (valid_i_gather_nw[5][22]),
    .data_o_gather_nw               (data_i_gather_nw[5][22]),
    .ready_i_gather_nw              (ready_o_gather_nw[5][22]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[5][22]),
    .data_i_merge_nw                (data_o_merge_nw[5][22]),
    .ready_o_merge_nw               (ready_i_merge_nw[5][22]),
    .valid_o_merge_nw               (valid_i_merge_nw[5][22]),
    .data_o_merge_nw                (data_i_merge_nw[5][22]),
    .ready_i_merge_nw               (ready_o_merge_nw[5][22]),

    .valid_i_cast_pe                (cast_valid_i_5_22),
    .data_i_cast_pe                 (cast_data_i_5_22),
    .ready_o_cast_pe                (cast_ready_o_5_22),
    .valid_o_cast_pe                (cast_valid_o_5_22),
    .data_o_cast_pe                 (cast_data_o_5_22),
    .ready_i_cast_pe                (cast_ready_i_5_22),

    .valid_i_merge_pe               (merge_valid_i_5_22),
    .data_i_merge_pe                (merge_data_i_5_22),
    .ready_o_merge_pe               (merge_ready_o_5_22),
    .valid_o_merge_pe               (merge_valid_o_5_22),
    .data_o_merge_pe                (merge_data_o_5_22),
    .ready_i_merge_pe               (merge_ready_i_5_22),

    .valid_i_gather_pe              (gather_valid_i_5_22),
    .data_i_gather_pe               (gather_data_i_5_22),
    .ready_o_gather_pe              (gather_ready_o_5_22),
    .valid_o_gather_pe              (gather_valid_o_5_22),
    .data_o_gather_pe               (gather_data_o_5_22),
    .ready_i_gather_pe              (gather_ready_i_5_22),

    .credit_upd                     (credit_upd[5][22])
);


network_interface #(
    .cast_out                       (cast_out_5_23),
    .gather_out                     (gather_out_5_23),
    .cast_sid                       (cast_sid_5_23),
    .gather_sid                     (gather_sid_5_23)
)ni_5_23(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[5][23]),
    .data_i_cast_nw                 (data_o_cast_nw[5][23]),
    .ready_o_cast_nw                (ready_i_cast_nw[5][23]),
    .valid_o_cast_nw                (valid_i_cast_nw[5][23]),
    .data_o_cast_nw                 (data_i_cast_nw[5][23]),
    .ready_i_cast_nw                (ready_o_cast_nw[5][23]),

    .valid_i_gather_nw              (valid_o_gather_nw[5][23]),
    .data_i_gather_nw               (data_o_gather_nw[5][23]),
    .ready_o_gather_nw              (ready_i_gather_nw[5][23]),
    .valid_o_gather_nw              (valid_i_gather_nw[5][23]),
    .data_o_gather_nw               (data_i_gather_nw[5][23]),
    .ready_i_gather_nw              (ready_o_gather_nw[5][23]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[5][23]),
    .data_i_merge_nw                (data_o_merge_nw[5][23]),
    .ready_o_merge_nw               (ready_i_merge_nw[5][23]),
    .valid_o_merge_nw               (valid_i_merge_nw[5][23]),
    .data_o_merge_nw                (data_i_merge_nw[5][23]),
    .ready_i_merge_nw               (ready_o_merge_nw[5][23]),

    .valid_i_cast_pe                (cast_valid_i_5_23),
    .data_i_cast_pe                 (cast_data_i_5_23),
    .ready_o_cast_pe                (cast_ready_o_5_23),
    .valid_o_cast_pe                (cast_valid_o_5_23),
    .data_o_cast_pe                 (cast_data_o_5_23),
    .ready_i_cast_pe                (cast_ready_i_5_23),

    .valid_i_merge_pe               (merge_valid_i_5_23),
    .data_i_merge_pe                (merge_data_i_5_23),
    .ready_o_merge_pe               (merge_ready_o_5_23),
    .valid_o_merge_pe               (merge_valid_o_5_23),
    .data_o_merge_pe                (merge_data_o_5_23),
    .ready_i_merge_pe               (merge_ready_i_5_23),

    .valid_i_gather_pe              (gather_valid_i_5_23),
    .data_i_gather_pe               (gather_data_i_5_23),
    .ready_o_gather_pe              (gather_ready_o_5_23),
    .valid_o_gather_pe              (gather_valid_o_5_23),
    .data_o_gather_pe               (gather_data_o_5_23),
    .ready_i_gather_pe              (gather_ready_i_5_23),

    .credit_upd                     (credit_upd[5][23])
);


network_interface #(
    .cast_out                       (cast_out_5_24),
    .gather_out                     (gather_out_5_24),
    .cast_sid                       (cast_sid_5_24),
    .gather_sid                     (gather_sid_5_24)
)ni_5_24(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[5][24]),
    .data_i_cast_nw                 (data_o_cast_nw[5][24]),
    .ready_o_cast_nw                (ready_i_cast_nw[5][24]),
    .valid_o_cast_nw                (valid_i_cast_nw[5][24]),
    .data_o_cast_nw                 (data_i_cast_nw[5][24]),
    .ready_i_cast_nw                (ready_o_cast_nw[5][24]),

    .valid_i_gather_nw              (valid_o_gather_nw[5][24]),
    .data_i_gather_nw               (data_o_gather_nw[5][24]),
    .ready_o_gather_nw              (ready_i_gather_nw[5][24]),
    .valid_o_gather_nw              (valid_i_gather_nw[5][24]),
    .data_o_gather_nw               (data_i_gather_nw[5][24]),
    .ready_i_gather_nw              (ready_o_gather_nw[5][24]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[5][24]),
    .data_i_merge_nw                (data_o_merge_nw[5][24]),
    .ready_o_merge_nw               (ready_i_merge_nw[5][24]),
    .valid_o_merge_nw               (valid_i_merge_nw[5][24]),
    .data_o_merge_nw                (data_i_merge_nw[5][24]),
    .ready_i_merge_nw               (ready_o_merge_nw[5][24]),

    .valid_i_cast_pe                (cast_valid_i_5_24),
    .data_i_cast_pe                 (cast_data_i_5_24),
    .ready_o_cast_pe                (cast_ready_o_5_24),
    .valid_o_cast_pe                (cast_valid_o_5_24),
    .data_o_cast_pe                 (cast_data_o_5_24),
    .ready_i_cast_pe                (cast_ready_i_5_24),

    .valid_i_merge_pe               (merge_valid_i_5_24),
    .data_i_merge_pe                (merge_data_i_5_24),
    .ready_o_merge_pe               (merge_ready_o_5_24),
    .valid_o_merge_pe               (merge_valid_o_5_24),
    .data_o_merge_pe                (merge_data_o_5_24),
    .ready_i_merge_pe               (merge_ready_i_5_24),

    .valid_i_gather_pe              (gather_valid_i_5_24),
    .data_i_gather_pe               (gather_data_i_5_24),
    .ready_o_gather_pe              (gather_ready_o_5_24),
    .valid_o_gather_pe              (gather_valid_o_5_24),
    .data_o_gather_pe               (gather_data_o_5_24),
    .ready_i_gather_pe              (gather_ready_i_5_24),

    .credit_upd                     (credit_upd[5][24])
);


network_interface #(
    .cast_out                       (cast_out_6_0),
    .gather_out                     (gather_out_6_0),
    .cast_sid                       (cast_sid_6_0),
    .gather_sid                     (gather_sid_6_0)
)ni_6_0(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[6][0]),
    .data_i_cast_nw                 (data_o_cast_nw[6][0]),
    .ready_o_cast_nw                (ready_i_cast_nw[6][0]),
    .valid_o_cast_nw                (valid_i_cast_nw[6][0]),
    .data_o_cast_nw                 (data_i_cast_nw[6][0]),
    .ready_i_cast_nw                (ready_o_cast_nw[6][0]),

    .valid_i_gather_nw              (valid_o_gather_nw[6][0]),
    .data_i_gather_nw               (data_o_gather_nw[6][0]),
    .ready_o_gather_nw              (ready_i_gather_nw[6][0]),
    .valid_o_gather_nw              (valid_i_gather_nw[6][0]),
    .data_o_gather_nw               (data_i_gather_nw[6][0]),
    .ready_i_gather_nw              (ready_o_gather_nw[6][0]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[6][0]),
    .data_i_merge_nw                (data_o_merge_nw[6][0]),
    .ready_o_merge_nw               (ready_i_merge_nw[6][0]),
    .valid_o_merge_nw               (valid_i_merge_nw[6][0]),
    .data_o_merge_nw                (data_i_merge_nw[6][0]),
    .ready_i_merge_nw               (ready_o_merge_nw[6][0]),

    .valid_i_cast_pe                (cast_valid_i_6_0),
    .data_i_cast_pe                 (cast_data_i_6_0),
    .ready_o_cast_pe                (cast_ready_o_6_0),
    .valid_o_cast_pe                (cast_valid_o_6_0),
    .data_o_cast_pe                 (cast_data_o_6_0),
    .ready_i_cast_pe                (cast_ready_i_6_0),

    .valid_i_merge_pe               (merge_valid_i_6_0),
    .data_i_merge_pe                (merge_data_i_6_0),
    .ready_o_merge_pe               (merge_ready_o_6_0),
    .valid_o_merge_pe               (merge_valid_o_6_0),
    .data_o_merge_pe                (merge_data_o_6_0),
    .ready_i_merge_pe               (merge_ready_i_6_0),

    .valid_i_gather_pe              (gather_valid_i_6_0),
    .data_i_gather_pe               (gather_data_i_6_0),
    .ready_o_gather_pe              (gather_ready_o_6_0),
    .valid_o_gather_pe              (gather_valid_o_6_0),
    .data_o_gather_pe               (gather_data_o_6_0),
    .ready_i_gather_pe              (gather_ready_i_6_0),

    .credit_upd                     (credit_upd[6][0])
);


network_interface #(
    .cast_out                       (cast_out_6_1),
    .gather_out                     (gather_out_6_1),
    .cast_sid                       (cast_sid_6_1),
    .gather_sid                     (gather_sid_6_1)
)ni_6_1(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[6][1]),
    .data_i_cast_nw                 (data_o_cast_nw[6][1]),
    .ready_o_cast_nw                (ready_i_cast_nw[6][1]),
    .valid_o_cast_nw                (valid_i_cast_nw[6][1]),
    .data_o_cast_nw                 (data_i_cast_nw[6][1]),
    .ready_i_cast_nw                (ready_o_cast_nw[6][1]),

    .valid_i_gather_nw              (valid_o_gather_nw[6][1]),
    .data_i_gather_nw               (data_o_gather_nw[6][1]),
    .ready_o_gather_nw              (ready_i_gather_nw[6][1]),
    .valid_o_gather_nw              (valid_i_gather_nw[6][1]),
    .data_o_gather_nw               (data_i_gather_nw[6][1]),
    .ready_i_gather_nw              (ready_o_gather_nw[6][1]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[6][1]),
    .data_i_merge_nw                (data_o_merge_nw[6][1]),
    .ready_o_merge_nw               (ready_i_merge_nw[6][1]),
    .valid_o_merge_nw               (valid_i_merge_nw[6][1]),
    .data_o_merge_nw                (data_i_merge_nw[6][1]),
    .ready_i_merge_nw               (ready_o_merge_nw[6][1]),

    .valid_i_cast_pe                (cast_valid_i_6_1),
    .data_i_cast_pe                 (cast_data_i_6_1),
    .ready_o_cast_pe                (cast_ready_o_6_1),
    .valid_o_cast_pe                (cast_valid_o_6_1),
    .data_o_cast_pe                 (cast_data_o_6_1),
    .ready_i_cast_pe                (cast_ready_i_6_1),

    .valid_i_merge_pe               (merge_valid_i_6_1),
    .data_i_merge_pe                (merge_data_i_6_1),
    .ready_o_merge_pe               (merge_ready_o_6_1),
    .valid_o_merge_pe               (merge_valid_o_6_1),
    .data_o_merge_pe                (merge_data_o_6_1),
    .ready_i_merge_pe               (merge_ready_i_6_1),

    .valid_i_gather_pe              (gather_valid_i_6_1),
    .data_i_gather_pe               (gather_data_i_6_1),
    .ready_o_gather_pe              (gather_ready_o_6_1),
    .valid_o_gather_pe              (gather_valid_o_6_1),
    .data_o_gather_pe               (gather_data_o_6_1),
    .ready_i_gather_pe              (gather_ready_i_6_1),

    .credit_upd                     (credit_upd[6][1])
);


network_interface #(
    .cast_out                       (cast_out_6_2),
    .gather_out                     (gather_out_6_2),
    .cast_sid                       (cast_sid_6_2),
    .gather_sid                     (gather_sid_6_2)
)ni_6_2(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[6][2]),
    .data_i_cast_nw                 (data_o_cast_nw[6][2]),
    .ready_o_cast_nw                (ready_i_cast_nw[6][2]),
    .valid_o_cast_nw                (valid_i_cast_nw[6][2]),
    .data_o_cast_nw                 (data_i_cast_nw[6][2]),
    .ready_i_cast_nw                (ready_o_cast_nw[6][2]),

    .valid_i_gather_nw              (valid_o_gather_nw[6][2]),
    .data_i_gather_nw               (data_o_gather_nw[6][2]),
    .ready_o_gather_nw              (ready_i_gather_nw[6][2]),
    .valid_o_gather_nw              (valid_i_gather_nw[6][2]),
    .data_o_gather_nw               (data_i_gather_nw[6][2]),
    .ready_i_gather_nw              (ready_o_gather_nw[6][2]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[6][2]),
    .data_i_merge_nw                (data_o_merge_nw[6][2]),
    .ready_o_merge_nw               (ready_i_merge_nw[6][2]),
    .valid_o_merge_nw               (valid_i_merge_nw[6][2]),
    .data_o_merge_nw                (data_i_merge_nw[6][2]),
    .ready_i_merge_nw               (ready_o_merge_nw[6][2]),

    .valid_i_cast_pe                (cast_valid_i_6_2),
    .data_i_cast_pe                 (cast_data_i_6_2),
    .ready_o_cast_pe                (cast_ready_o_6_2),
    .valid_o_cast_pe                (cast_valid_o_6_2),
    .data_o_cast_pe                 (cast_data_o_6_2),
    .ready_i_cast_pe                (cast_ready_i_6_2),

    .valid_i_merge_pe               (merge_valid_i_6_2),
    .data_i_merge_pe                (merge_data_i_6_2),
    .ready_o_merge_pe               (merge_ready_o_6_2),
    .valid_o_merge_pe               (merge_valid_o_6_2),
    .data_o_merge_pe                (merge_data_o_6_2),
    .ready_i_merge_pe               (merge_ready_i_6_2),

    .valid_i_gather_pe              (gather_valid_i_6_2),
    .data_i_gather_pe               (gather_data_i_6_2),
    .ready_o_gather_pe              (gather_ready_o_6_2),
    .valid_o_gather_pe              (gather_valid_o_6_2),
    .data_o_gather_pe               (gather_data_o_6_2),
    .ready_i_gather_pe              (gather_ready_i_6_2),

    .credit_upd                     (credit_upd[6][2])
);


network_interface #(
    .cast_out                       (cast_out_6_3),
    .gather_out                     (gather_out_6_3),
    .cast_sid                       (cast_sid_6_3),
    .gather_sid                     (gather_sid_6_3)
)ni_6_3(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[6][3]),
    .data_i_cast_nw                 (data_o_cast_nw[6][3]),
    .ready_o_cast_nw                (ready_i_cast_nw[6][3]),
    .valid_o_cast_nw                (valid_i_cast_nw[6][3]),
    .data_o_cast_nw                 (data_i_cast_nw[6][3]),
    .ready_i_cast_nw                (ready_o_cast_nw[6][3]),

    .valid_i_gather_nw              (valid_o_gather_nw[6][3]),
    .data_i_gather_nw               (data_o_gather_nw[6][3]),
    .ready_o_gather_nw              (ready_i_gather_nw[6][3]),
    .valid_o_gather_nw              (valid_i_gather_nw[6][3]),
    .data_o_gather_nw               (data_i_gather_nw[6][3]),
    .ready_i_gather_nw              (ready_o_gather_nw[6][3]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[6][3]),
    .data_i_merge_nw                (data_o_merge_nw[6][3]),
    .ready_o_merge_nw               (ready_i_merge_nw[6][3]),
    .valid_o_merge_nw               (valid_i_merge_nw[6][3]),
    .data_o_merge_nw                (data_i_merge_nw[6][3]),
    .ready_i_merge_nw               (ready_o_merge_nw[6][3]),

    .valid_i_cast_pe                (cast_valid_i_6_3),
    .data_i_cast_pe                 (cast_data_i_6_3),
    .ready_o_cast_pe                (cast_ready_o_6_3),
    .valid_o_cast_pe                (cast_valid_o_6_3),
    .data_o_cast_pe                 (cast_data_o_6_3),
    .ready_i_cast_pe                (cast_ready_i_6_3),

    .valid_i_merge_pe               (merge_valid_i_6_3),
    .data_i_merge_pe                (merge_data_i_6_3),
    .ready_o_merge_pe               (merge_ready_o_6_3),
    .valid_o_merge_pe               (merge_valid_o_6_3),
    .data_o_merge_pe                (merge_data_o_6_3),
    .ready_i_merge_pe               (merge_ready_i_6_3),

    .valid_i_gather_pe              (gather_valid_i_6_3),
    .data_i_gather_pe               (gather_data_i_6_3),
    .ready_o_gather_pe              (gather_ready_o_6_3),
    .valid_o_gather_pe              (gather_valid_o_6_3),
    .data_o_gather_pe               (gather_data_o_6_3),
    .ready_i_gather_pe              (gather_ready_i_6_3),

    .credit_upd                     (credit_upd[6][3])
);


network_interface #(
    .cast_out                       (cast_out_6_4),
    .gather_out                     (gather_out_6_4),
    .cast_sid                       (cast_sid_6_4),
    .gather_sid                     (gather_sid_6_4)
)ni_6_4(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[6][4]),
    .data_i_cast_nw                 (data_o_cast_nw[6][4]),
    .ready_o_cast_nw                (ready_i_cast_nw[6][4]),
    .valid_o_cast_nw                (valid_i_cast_nw[6][4]),
    .data_o_cast_nw                 (data_i_cast_nw[6][4]),
    .ready_i_cast_nw                (ready_o_cast_nw[6][4]),

    .valid_i_gather_nw              (valid_o_gather_nw[6][4]),
    .data_i_gather_nw               (data_o_gather_nw[6][4]),
    .ready_o_gather_nw              (ready_i_gather_nw[6][4]),
    .valid_o_gather_nw              (valid_i_gather_nw[6][4]),
    .data_o_gather_nw               (data_i_gather_nw[6][4]),
    .ready_i_gather_nw              (ready_o_gather_nw[6][4]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[6][4]),
    .data_i_merge_nw                (data_o_merge_nw[6][4]),
    .ready_o_merge_nw               (ready_i_merge_nw[6][4]),
    .valid_o_merge_nw               (valid_i_merge_nw[6][4]),
    .data_o_merge_nw                (data_i_merge_nw[6][4]),
    .ready_i_merge_nw               (ready_o_merge_nw[6][4]),

    .valid_i_cast_pe                (cast_valid_i_6_4),
    .data_i_cast_pe                 (cast_data_i_6_4),
    .ready_o_cast_pe                (cast_ready_o_6_4),
    .valid_o_cast_pe                (cast_valid_o_6_4),
    .data_o_cast_pe                 (cast_data_o_6_4),
    .ready_i_cast_pe                (cast_ready_i_6_4),

    .valid_i_merge_pe               (merge_valid_i_6_4),
    .data_i_merge_pe                (merge_data_i_6_4),
    .ready_o_merge_pe               (merge_ready_o_6_4),
    .valid_o_merge_pe               (merge_valid_o_6_4),
    .data_o_merge_pe                (merge_data_o_6_4),
    .ready_i_merge_pe               (merge_ready_i_6_4),

    .valid_i_gather_pe              (gather_valid_i_6_4),
    .data_i_gather_pe               (gather_data_i_6_4),
    .ready_o_gather_pe              (gather_ready_o_6_4),
    .valid_o_gather_pe              (gather_valid_o_6_4),
    .data_o_gather_pe               (gather_data_o_6_4),
    .ready_i_gather_pe              (gather_ready_i_6_4),

    .credit_upd                     (credit_upd[6][4])
);


network_interface #(
    .cast_out                       (cast_out_6_5),
    .gather_out                     (gather_out_6_5),
    .cast_sid                       (cast_sid_6_5),
    .gather_sid                     (gather_sid_6_5)
)ni_6_5(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[6][5]),
    .data_i_cast_nw                 (data_o_cast_nw[6][5]),
    .ready_o_cast_nw                (ready_i_cast_nw[6][5]),
    .valid_o_cast_nw                (valid_i_cast_nw[6][5]),
    .data_o_cast_nw                 (data_i_cast_nw[6][5]),
    .ready_i_cast_nw                (ready_o_cast_nw[6][5]),

    .valid_i_gather_nw              (valid_o_gather_nw[6][5]),
    .data_i_gather_nw               (data_o_gather_nw[6][5]),
    .ready_o_gather_nw              (ready_i_gather_nw[6][5]),
    .valid_o_gather_nw              (valid_i_gather_nw[6][5]),
    .data_o_gather_nw               (data_i_gather_nw[6][5]),
    .ready_i_gather_nw              (ready_o_gather_nw[6][5]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[6][5]),
    .data_i_merge_nw                (data_o_merge_nw[6][5]),
    .ready_o_merge_nw               (ready_i_merge_nw[6][5]),
    .valid_o_merge_nw               (valid_i_merge_nw[6][5]),
    .data_o_merge_nw                (data_i_merge_nw[6][5]),
    .ready_i_merge_nw               (ready_o_merge_nw[6][5]),

    .valid_i_cast_pe                (cast_valid_i_6_5),
    .data_i_cast_pe                 (cast_data_i_6_5),
    .ready_o_cast_pe                (cast_ready_o_6_5),
    .valid_o_cast_pe                (cast_valid_o_6_5),
    .data_o_cast_pe                 (cast_data_o_6_5),
    .ready_i_cast_pe                (cast_ready_i_6_5),

    .valid_i_merge_pe               (merge_valid_i_6_5),
    .data_i_merge_pe                (merge_data_i_6_5),
    .ready_o_merge_pe               (merge_ready_o_6_5),
    .valid_o_merge_pe               (merge_valid_o_6_5),
    .data_o_merge_pe                (merge_data_o_6_5),
    .ready_i_merge_pe               (merge_ready_i_6_5),

    .valid_i_gather_pe              (gather_valid_i_6_5),
    .data_i_gather_pe               (gather_data_i_6_5),
    .ready_o_gather_pe              (gather_ready_o_6_5),
    .valid_o_gather_pe              (gather_valid_o_6_5),
    .data_o_gather_pe               (gather_data_o_6_5),
    .ready_i_gather_pe              (gather_ready_i_6_5),

    .credit_upd                     (credit_upd[6][5])
);


network_interface #(
    .cast_out                       (cast_out_6_6),
    .gather_out                     (gather_out_6_6),
    .cast_sid                       (cast_sid_6_6),
    .gather_sid                     (gather_sid_6_6)
)ni_6_6(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[6][6]),
    .data_i_cast_nw                 (data_o_cast_nw[6][6]),
    .ready_o_cast_nw                (ready_i_cast_nw[6][6]),
    .valid_o_cast_nw                (valid_i_cast_nw[6][6]),
    .data_o_cast_nw                 (data_i_cast_nw[6][6]),
    .ready_i_cast_nw                (ready_o_cast_nw[6][6]),

    .valid_i_gather_nw              (valid_o_gather_nw[6][6]),
    .data_i_gather_nw               (data_o_gather_nw[6][6]),
    .ready_o_gather_nw              (ready_i_gather_nw[6][6]),
    .valid_o_gather_nw              (valid_i_gather_nw[6][6]),
    .data_o_gather_nw               (data_i_gather_nw[6][6]),
    .ready_i_gather_nw              (ready_o_gather_nw[6][6]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[6][6]),
    .data_i_merge_nw                (data_o_merge_nw[6][6]),
    .ready_o_merge_nw               (ready_i_merge_nw[6][6]),
    .valid_o_merge_nw               (valid_i_merge_nw[6][6]),
    .data_o_merge_nw                (data_i_merge_nw[6][6]),
    .ready_i_merge_nw               (ready_o_merge_nw[6][6]),

    .valid_i_cast_pe                (cast_valid_i_6_6),
    .data_i_cast_pe                 (cast_data_i_6_6),
    .ready_o_cast_pe                (cast_ready_o_6_6),
    .valid_o_cast_pe                (cast_valid_o_6_6),
    .data_o_cast_pe                 (cast_data_o_6_6),
    .ready_i_cast_pe                (cast_ready_i_6_6),

    .valid_i_merge_pe               (merge_valid_i_6_6),
    .data_i_merge_pe                (merge_data_i_6_6),
    .ready_o_merge_pe               (merge_ready_o_6_6),
    .valid_o_merge_pe               (merge_valid_o_6_6),
    .data_o_merge_pe                (merge_data_o_6_6),
    .ready_i_merge_pe               (merge_ready_i_6_6),

    .valid_i_gather_pe              (gather_valid_i_6_6),
    .data_i_gather_pe               (gather_data_i_6_6),
    .ready_o_gather_pe              (gather_ready_o_6_6),
    .valid_o_gather_pe              (gather_valid_o_6_6),
    .data_o_gather_pe               (gather_data_o_6_6),
    .ready_i_gather_pe              (gather_ready_i_6_6),

    .credit_upd                     (credit_upd[6][6])
);


network_interface #(
    .cast_out                       (cast_out_6_7),
    .gather_out                     (gather_out_6_7),
    .cast_sid                       (cast_sid_6_7),
    .gather_sid                     (gather_sid_6_7)
)ni_6_7(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[6][7]),
    .data_i_cast_nw                 (data_o_cast_nw[6][7]),
    .ready_o_cast_nw                (ready_i_cast_nw[6][7]),
    .valid_o_cast_nw                (valid_i_cast_nw[6][7]),
    .data_o_cast_nw                 (data_i_cast_nw[6][7]),
    .ready_i_cast_nw                (ready_o_cast_nw[6][7]),

    .valid_i_gather_nw              (valid_o_gather_nw[6][7]),
    .data_i_gather_nw               (data_o_gather_nw[6][7]),
    .ready_o_gather_nw              (ready_i_gather_nw[6][7]),
    .valid_o_gather_nw              (valid_i_gather_nw[6][7]),
    .data_o_gather_nw               (data_i_gather_nw[6][7]),
    .ready_i_gather_nw              (ready_o_gather_nw[6][7]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[6][7]),
    .data_i_merge_nw                (data_o_merge_nw[6][7]),
    .ready_o_merge_nw               (ready_i_merge_nw[6][7]),
    .valid_o_merge_nw               (valid_i_merge_nw[6][7]),
    .data_o_merge_nw                (data_i_merge_nw[6][7]),
    .ready_i_merge_nw               (ready_o_merge_nw[6][7]),

    .valid_i_cast_pe                (cast_valid_i_6_7),
    .data_i_cast_pe                 (cast_data_i_6_7),
    .ready_o_cast_pe                (cast_ready_o_6_7),
    .valid_o_cast_pe                (cast_valid_o_6_7),
    .data_o_cast_pe                 (cast_data_o_6_7),
    .ready_i_cast_pe                (cast_ready_i_6_7),

    .valid_i_merge_pe               (merge_valid_i_6_7),
    .data_i_merge_pe                (merge_data_i_6_7),
    .ready_o_merge_pe               (merge_ready_o_6_7),
    .valid_o_merge_pe               (merge_valid_o_6_7),
    .data_o_merge_pe                (merge_data_o_6_7),
    .ready_i_merge_pe               (merge_ready_i_6_7),

    .valid_i_gather_pe              (gather_valid_i_6_7),
    .data_i_gather_pe               (gather_data_i_6_7),
    .ready_o_gather_pe              (gather_ready_o_6_7),
    .valid_o_gather_pe              (gather_valid_o_6_7),
    .data_o_gather_pe               (gather_data_o_6_7),
    .ready_i_gather_pe              (gather_ready_i_6_7),

    .credit_upd                     (credit_upd[6][7])
);


network_interface #(
    .cast_out                       (cast_out_6_8),
    .gather_out                     (gather_out_6_8),
    .cast_sid                       (cast_sid_6_8),
    .gather_sid                     (gather_sid_6_8)
)ni_6_8(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[6][8]),
    .data_i_cast_nw                 (data_o_cast_nw[6][8]),
    .ready_o_cast_nw                (ready_i_cast_nw[6][8]),
    .valid_o_cast_nw                (valid_i_cast_nw[6][8]),
    .data_o_cast_nw                 (data_i_cast_nw[6][8]),
    .ready_i_cast_nw                (ready_o_cast_nw[6][8]),

    .valid_i_gather_nw              (valid_o_gather_nw[6][8]),
    .data_i_gather_nw               (data_o_gather_nw[6][8]),
    .ready_o_gather_nw              (ready_i_gather_nw[6][8]),
    .valid_o_gather_nw              (valid_i_gather_nw[6][8]),
    .data_o_gather_nw               (data_i_gather_nw[6][8]),
    .ready_i_gather_nw              (ready_o_gather_nw[6][8]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[6][8]),
    .data_i_merge_nw                (data_o_merge_nw[6][8]),
    .ready_o_merge_nw               (ready_i_merge_nw[6][8]),
    .valid_o_merge_nw               (valid_i_merge_nw[6][8]),
    .data_o_merge_nw                (data_i_merge_nw[6][8]),
    .ready_i_merge_nw               (ready_o_merge_nw[6][8]),

    .valid_i_cast_pe                (cast_valid_i_6_8),
    .data_i_cast_pe                 (cast_data_i_6_8),
    .ready_o_cast_pe                (cast_ready_o_6_8),
    .valid_o_cast_pe                (cast_valid_o_6_8),
    .data_o_cast_pe                 (cast_data_o_6_8),
    .ready_i_cast_pe                (cast_ready_i_6_8),

    .valid_i_merge_pe               (merge_valid_i_6_8),
    .data_i_merge_pe                (merge_data_i_6_8),
    .ready_o_merge_pe               (merge_ready_o_6_8),
    .valid_o_merge_pe               (merge_valid_o_6_8),
    .data_o_merge_pe                (merge_data_o_6_8),
    .ready_i_merge_pe               (merge_ready_i_6_8),

    .valid_i_gather_pe              (gather_valid_i_6_8),
    .data_i_gather_pe               (gather_data_i_6_8),
    .ready_o_gather_pe              (gather_ready_o_6_8),
    .valid_o_gather_pe              (gather_valid_o_6_8),
    .data_o_gather_pe               (gather_data_o_6_8),
    .ready_i_gather_pe              (gather_ready_i_6_8),

    .credit_upd                     (credit_upd[6][8])
);


network_interface #(
    .cast_out                       (cast_out_6_9),
    .gather_out                     (gather_out_6_9),
    .cast_sid                       (cast_sid_6_9),
    .gather_sid                     (gather_sid_6_9)
)ni_6_9(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[6][9]),
    .data_i_cast_nw                 (data_o_cast_nw[6][9]),
    .ready_o_cast_nw                (ready_i_cast_nw[6][9]),
    .valid_o_cast_nw                (valid_i_cast_nw[6][9]),
    .data_o_cast_nw                 (data_i_cast_nw[6][9]),
    .ready_i_cast_nw                (ready_o_cast_nw[6][9]),

    .valid_i_gather_nw              (valid_o_gather_nw[6][9]),
    .data_i_gather_nw               (data_o_gather_nw[6][9]),
    .ready_o_gather_nw              (ready_i_gather_nw[6][9]),
    .valid_o_gather_nw              (valid_i_gather_nw[6][9]),
    .data_o_gather_nw               (data_i_gather_nw[6][9]),
    .ready_i_gather_nw              (ready_o_gather_nw[6][9]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[6][9]),
    .data_i_merge_nw                (data_o_merge_nw[6][9]),
    .ready_o_merge_nw               (ready_i_merge_nw[6][9]),
    .valid_o_merge_nw               (valid_i_merge_nw[6][9]),
    .data_o_merge_nw                (data_i_merge_nw[6][9]),
    .ready_i_merge_nw               (ready_o_merge_nw[6][9]),

    .valid_i_cast_pe                (cast_valid_i_6_9),
    .data_i_cast_pe                 (cast_data_i_6_9),
    .ready_o_cast_pe                (cast_ready_o_6_9),
    .valid_o_cast_pe                (cast_valid_o_6_9),
    .data_o_cast_pe                 (cast_data_o_6_9),
    .ready_i_cast_pe                (cast_ready_i_6_9),

    .valid_i_merge_pe               (merge_valid_i_6_9),
    .data_i_merge_pe                (merge_data_i_6_9),
    .ready_o_merge_pe               (merge_ready_o_6_9),
    .valid_o_merge_pe               (merge_valid_o_6_9),
    .data_o_merge_pe                (merge_data_o_6_9),
    .ready_i_merge_pe               (merge_ready_i_6_9),

    .valid_i_gather_pe              (gather_valid_i_6_9),
    .data_i_gather_pe               (gather_data_i_6_9),
    .ready_o_gather_pe              (gather_ready_o_6_9),
    .valid_o_gather_pe              (gather_valid_o_6_9),
    .data_o_gather_pe               (gather_data_o_6_9),
    .ready_i_gather_pe              (gather_ready_i_6_9),

    .credit_upd                     (credit_upd[6][9])
);


network_interface #(
    .cast_out                       (cast_out_6_10),
    .gather_out                     (gather_out_6_10),
    .cast_sid                       (cast_sid_6_10),
    .gather_sid                     (gather_sid_6_10)
)ni_6_10(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[6][10]),
    .data_i_cast_nw                 (data_o_cast_nw[6][10]),
    .ready_o_cast_nw                (ready_i_cast_nw[6][10]),
    .valid_o_cast_nw                (valid_i_cast_nw[6][10]),
    .data_o_cast_nw                 (data_i_cast_nw[6][10]),
    .ready_i_cast_nw                (ready_o_cast_nw[6][10]),

    .valid_i_gather_nw              (valid_o_gather_nw[6][10]),
    .data_i_gather_nw               (data_o_gather_nw[6][10]),
    .ready_o_gather_nw              (ready_i_gather_nw[6][10]),
    .valid_o_gather_nw              (valid_i_gather_nw[6][10]),
    .data_o_gather_nw               (data_i_gather_nw[6][10]),
    .ready_i_gather_nw              (ready_o_gather_nw[6][10]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[6][10]),
    .data_i_merge_nw                (data_o_merge_nw[6][10]),
    .ready_o_merge_nw               (ready_i_merge_nw[6][10]),
    .valid_o_merge_nw               (valid_i_merge_nw[6][10]),
    .data_o_merge_nw                (data_i_merge_nw[6][10]),
    .ready_i_merge_nw               (ready_o_merge_nw[6][10]),

    .valid_i_cast_pe                (cast_valid_i_6_10),
    .data_i_cast_pe                 (cast_data_i_6_10),
    .ready_o_cast_pe                (cast_ready_o_6_10),
    .valid_o_cast_pe                (cast_valid_o_6_10),
    .data_o_cast_pe                 (cast_data_o_6_10),
    .ready_i_cast_pe                (cast_ready_i_6_10),

    .valid_i_merge_pe               (merge_valid_i_6_10),
    .data_i_merge_pe                (merge_data_i_6_10),
    .ready_o_merge_pe               (merge_ready_o_6_10),
    .valid_o_merge_pe               (merge_valid_o_6_10),
    .data_o_merge_pe                (merge_data_o_6_10),
    .ready_i_merge_pe               (merge_ready_i_6_10),

    .valid_i_gather_pe              (gather_valid_i_6_10),
    .data_i_gather_pe               (gather_data_i_6_10),
    .ready_o_gather_pe              (gather_ready_o_6_10),
    .valid_o_gather_pe              (gather_valid_o_6_10),
    .data_o_gather_pe               (gather_data_o_6_10),
    .ready_i_gather_pe              (gather_ready_i_6_10),

    .credit_upd                     (credit_upd[6][10])
);


network_interface #(
    .cast_out                       (cast_out_6_11),
    .gather_out                     (gather_out_6_11),
    .cast_sid                       (cast_sid_6_11),
    .gather_sid                     (gather_sid_6_11)
)ni_6_11(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[6][11]),
    .data_i_cast_nw                 (data_o_cast_nw[6][11]),
    .ready_o_cast_nw                (ready_i_cast_nw[6][11]),
    .valid_o_cast_nw                (valid_i_cast_nw[6][11]),
    .data_o_cast_nw                 (data_i_cast_nw[6][11]),
    .ready_i_cast_nw                (ready_o_cast_nw[6][11]),

    .valid_i_gather_nw              (valid_o_gather_nw[6][11]),
    .data_i_gather_nw               (data_o_gather_nw[6][11]),
    .ready_o_gather_nw              (ready_i_gather_nw[6][11]),
    .valid_o_gather_nw              (valid_i_gather_nw[6][11]),
    .data_o_gather_nw               (data_i_gather_nw[6][11]),
    .ready_i_gather_nw              (ready_o_gather_nw[6][11]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[6][11]),
    .data_i_merge_nw                (data_o_merge_nw[6][11]),
    .ready_o_merge_nw               (ready_i_merge_nw[6][11]),
    .valid_o_merge_nw               (valid_i_merge_nw[6][11]),
    .data_o_merge_nw                (data_i_merge_nw[6][11]),
    .ready_i_merge_nw               (ready_o_merge_nw[6][11]),

    .valid_i_cast_pe                (cast_valid_i_6_11),
    .data_i_cast_pe                 (cast_data_i_6_11),
    .ready_o_cast_pe                (cast_ready_o_6_11),
    .valid_o_cast_pe                (cast_valid_o_6_11),
    .data_o_cast_pe                 (cast_data_o_6_11),
    .ready_i_cast_pe                (cast_ready_i_6_11),

    .valid_i_merge_pe               (merge_valid_i_6_11),
    .data_i_merge_pe                (merge_data_i_6_11),
    .ready_o_merge_pe               (merge_ready_o_6_11),
    .valid_o_merge_pe               (merge_valid_o_6_11),
    .data_o_merge_pe                (merge_data_o_6_11),
    .ready_i_merge_pe               (merge_ready_i_6_11),

    .valid_i_gather_pe              (gather_valid_i_6_11),
    .data_i_gather_pe               (gather_data_i_6_11),
    .ready_o_gather_pe              (gather_ready_o_6_11),
    .valid_o_gather_pe              (gather_valid_o_6_11),
    .data_o_gather_pe               (gather_data_o_6_11),
    .ready_i_gather_pe              (gather_ready_i_6_11),

    .credit_upd                     (credit_upd[6][11])
);


network_interface #(
    .cast_out                       (cast_out_6_12),
    .gather_out                     (gather_out_6_12),
    .cast_sid                       (cast_sid_6_12),
    .gather_sid                     (gather_sid_6_12)
)ni_6_12(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[6][12]),
    .data_i_cast_nw                 (data_o_cast_nw[6][12]),
    .ready_o_cast_nw                (ready_i_cast_nw[6][12]),
    .valid_o_cast_nw                (valid_i_cast_nw[6][12]),
    .data_o_cast_nw                 (data_i_cast_nw[6][12]),
    .ready_i_cast_nw                (ready_o_cast_nw[6][12]),

    .valid_i_gather_nw              (valid_o_gather_nw[6][12]),
    .data_i_gather_nw               (data_o_gather_nw[6][12]),
    .ready_o_gather_nw              (ready_i_gather_nw[6][12]),
    .valid_o_gather_nw              (valid_i_gather_nw[6][12]),
    .data_o_gather_nw               (data_i_gather_nw[6][12]),
    .ready_i_gather_nw              (ready_o_gather_nw[6][12]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[6][12]),
    .data_i_merge_nw                (data_o_merge_nw[6][12]),
    .ready_o_merge_nw               (ready_i_merge_nw[6][12]),
    .valid_o_merge_nw               (valid_i_merge_nw[6][12]),
    .data_o_merge_nw                (data_i_merge_nw[6][12]),
    .ready_i_merge_nw               (ready_o_merge_nw[6][12]),

    .valid_i_cast_pe                (cast_valid_i_6_12),
    .data_i_cast_pe                 (cast_data_i_6_12),
    .ready_o_cast_pe                (cast_ready_o_6_12),
    .valid_o_cast_pe                (cast_valid_o_6_12),
    .data_o_cast_pe                 (cast_data_o_6_12),
    .ready_i_cast_pe                (cast_ready_i_6_12),

    .valid_i_merge_pe               (merge_valid_i_6_12),
    .data_i_merge_pe                (merge_data_i_6_12),
    .ready_o_merge_pe               (merge_ready_o_6_12),
    .valid_o_merge_pe               (merge_valid_o_6_12),
    .data_o_merge_pe                (merge_data_o_6_12),
    .ready_i_merge_pe               (merge_ready_i_6_12),

    .valid_i_gather_pe              (gather_valid_i_6_12),
    .data_i_gather_pe               (gather_data_i_6_12),
    .ready_o_gather_pe              (gather_ready_o_6_12),
    .valid_o_gather_pe              (gather_valid_o_6_12),
    .data_o_gather_pe               (gather_data_o_6_12),
    .ready_i_gather_pe              (gather_ready_i_6_12),

    .credit_upd                     (credit_upd[6][12])
);


network_interface #(
    .cast_out                       (cast_out_6_13),
    .gather_out                     (gather_out_6_13),
    .cast_sid                       (cast_sid_6_13),
    .gather_sid                     (gather_sid_6_13)
)ni_6_13(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[6][13]),
    .data_i_cast_nw                 (data_o_cast_nw[6][13]),
    .ready_o_cast_nw                (ready_i_cast_nw[6][13]),
    .valid_o_cast_nw                (valid_i_cast_nw[6][13]),
    .data_o_cast_nw                 (data_i_cast_nw[6][13]),
    .ready_i_cast_nw                (ready_o_cast_nw[6][13]),

    .valid_i_gather_nw              (valid_o_gather_nw[6][13]),
    .data_i_gather_nw               (data_o_gather_nw[6][13]),
    .ready_o_gather_nw              (ready_i_gather_nw[6][13]),
    .valid_o_gather_nw              (valid_i_gather_nw[6][13]),
    .data_o_gather_nw               (data_i_gather_nw[6][13]),
    .ready_i_gather_nw              (ready_o_gather_nw[6][13]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[6][13]),
    .data_i_merge_nw                (data_o_merge_nw[6][13]),
    .ready_o_merge_nw               (ready_i_merge_nw[6][13]),
    .valid_o_merge_nw               (valid_i_merge_nw[6][13]),
    .data_o_merge_nw                (data_i_merge_nw[6][13]),
    .ready_i_merge_nw               (ready_o_merge_nw[6][13]),

    .valid_i_cast_pe                (cast_valid_i_6_13),
    .data_i_cast_pe                 (cast_data_i_6_13),
    .ready_o_cast_pe                (cast_ready_o_6_13),
    .valid_o_cast_pe                (cast_valid_o_6_13),
    .data_o_cast_pe                 (cast_data_o_6_13),
    .ready_i_cast_pe                (cast_ready_i_6_13),

    .valid_i_merge_pe               (merge_valid_i_6_13),
    .data_i_merge_pe                (merge_data_i_6_13),
    .ready_o_merge_pe               (merge_ready_o_6_13),
    .valid_o_merge_pe               (merge_valid_o_6_13),
    .data_o_merge_pe                (merge_data_o_6_13),
    .ready_i_merge_pe               (merge_ready_i_6_13),

    .valid_i_gather_pe              (gather_valid_i_6_13),
    .data_i_gather_pe               (gather_data_i_6_13),
    .ready_o_gather_pe              (gather_ready_o_6_13),
    .valid_o_gather_pe              (gather_valid_o_6_13),
    .data_o_gather_pe               (gather_data_o_6_13),
    .ready_i_gather_pe              (gather_ready_i_6_13),

    .credit_upd                     (credit_upd[6][13])
);


network_interface #(
    .cast_out                       (cast_out_6_14),
    .gather_out                     (gather_out_6_14),
    .cast_sid                       (cast_sid_6_14),
    .gather_sid                     (gather_sid_6_14)
)ni_6_14(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[6][14]),
    .data_i_cast_nw                 (data_o_cast_nw[6][14]),
    .ready_o_cast_nw                (ready_i_cast_nw[6][14]),
    .valid_o_cast_nw                (valid_i_cast_nw[6][14]),
    .data_o_cast_nw                 (data_i_cast_nw[6][14]),
    .ready_i_cast_nw                (ready_o_cast_nw[6][14]),

    .valid_i_gather_nw              (valid_o_gather_nw[6][14]),
    .data_i_gather_nw               (data_o_gather_nw[6][14]),
    .ready_o_gather_nw              (ready_i_gather_nw[6][14]),
    .valid_o_gather_nw              (valid_i_gather_nw[6][14]),
    .data_o_gather_nw               (data_i_gather_nw[6][14]),
    .ready_i_gather_nw              (ready_o_gather_nw[6][14]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[6][14]),
    .data_i_merge_nw                (data_o_merge_nw[6][14]),
    .ready_o_merge_nw               (ready_i_merge_nw[6][14]),
    .valid_o_merge_nw               (valid_i_merge_nw[6][14]),
    .data_o_merge_nw                (data_i_merge_nw[6][14]),
    .ready_i_merge_nw               (ready_o_merge_nw[6][14]),

    .valid_i_cast_pe                (cast_valid_i_6_14),
    .data_i_cast_pe                 (cast_data_i_6_14),
    .ready_o_cast_pe                (cast_ready_o_6_14),
    .valid_o_cast_pe                (cast_valid_o_6_14),
    .data_o_cast_pe                 (cast_data_o_6_14),
    .ready_i_cast_pe                (cast_ready_i_6_14),

    .valid_i_merge_pe               (merge_valid_i_6_14),
    .data_i_merge_pe                (merge_data_i_6_14),
    .ready_o_merge_pe               (merge_ready_o_6_14),
    .valid_o_merge_pe               (merge_valid_o_6_14),
    .data_o_merge_pe                (merge_data_o_6_14),
    .ready_i_merge_pe               (merge_ready_i_6_14),

    .valid_i_gather_pe              (gather_valid_i_6_14),
    .data_i_gather_pe               (gather_data_i_6_14),
    .ready_o_gather_pe              (gather_ready_o_6_14),
    .valid_o_gather_pe              (gather_valid_o_6_14),
    .data_o_gather_pe               (gather_data_o_6_14),
    .ready_i_gather_pe              (gather_ready_i_6_14),

    .credit_upd                     (credit_upd[6][14])
);


network_interface #(
    .cast_out                       (cast_out_6_15),
    .gather_out                     (gather_out_6_15),
    .cast_sid                       (cast_sid_6_15),
    .gather_sid                     (gather_sid_6_15)
)ni_6_15(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[6][15]),
    .data_i_cast_nw                 (data_o_cast_nw[6][15]),
    .ready_o_cast_nw                (ready_i_cast_nw[6][15]),
    .valid_o_cast_nw                (valid_i_cast_nw[6][15]),
    .data_o_cast_nw                 (data_i_cast_nw[6][15]),
    .ready_i_cast_nw                (ready_o_cast_nw[6][15]),

    .valid_i_gather_nw              (valid_o_gather_nw[6][15]),
    .data_i_gather_nw               (data_o_gather_nw[6][15]),
    .ready_o_gather_nw              (ready_i_gather_nw[6][15]),
    .valid_o_gather_nw              (valid_i_gather_nw[6][15]),
    .data_o_gather_nw               (data_i_gather_nw[6][15]),
    .ready_i_gather_nw              (ready_o_gather_nw[6][15]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[6][15]),
    .data_i_merge_nw                (data_o_merge_nw[6][15]),
    .ready_o_merge_nw               (ready_i_merge_nw[6][15]),
    .valid_o_merge_nw               (valid_i_merge_nw[6][15]),
    .data_o_merge_nw                (data_i_merge_nw[6][15]),
    .ready_i_merge_nw               (ready_o_merge_nw[6][15]),

    .valid_i_cast_pe                (cast_valid_i_6_15),
    .data_i_cast_pe                 (cast_data_i_6_15),
    .ready_o_cast_pe                (cast_ready_o_6_15),
    .valid_o_cast_pe                (cast_valid_o_6_15),
    .data_o_cast_pe                 (cast_data_o_6_15),
    .ready_i_cast_pe                (cast_ready_i_6_15),

    .valid_i_merge_pe               (merge_valid_i_6_15),
    .data_i_merge_pe                (merge_data_i_6_15),
    .ready_o_merge_pe               (merge_ready_o_6_15),
    .valid_o_merge_pe               (merge_valid_o_6_15),
    .data_o_merge_pe                (merge_data_o_6_15),
    .ready_i_merge_pe               (merge_ready_i_6_15),

    .valid_i_gather_pe              (gather_valid_i_6_15),
    .data_i_gather_pe               (gather_data_i_6_15),
    .ready_o_gather_pe              (gather_ready_o_6_15),
    .valid_o_gather_pe              (gather_valid_o_6_15),
    .data_o_gather_pe               (gather_data_o_6_15),
    .ready_i_gather_pe              (gather_ready_i_6_15),

    .credit_upd                     (credit_upd[6][15])
);


network_interface #(
    .cast_out                       (cast_out_6_16),
    .gather_out                     (gather_out_6_16),
    .cast_sid                       (cast_sid_6_16),
    .gather_sid                     (gather_sid_6_16)
)ni_6_16(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[6][16]),
    .data_i_cast_nw                 (data_o_cast_nw[6][16]),
    .ready_o_cast_nw                (ready_i_cast_nw[6][16]),
    .valid_o_cast_nw                (valid_i_cast_nw[6][16]),
    .data_o_cast_nw                 (data_i_cast_nw[6][16]),
    .ready_i_cast_nw                (ready_o_cast_nw[6][16]),

    .valid_i_gather_nw              (valid_o_gather_nw[6][16]),
    .data_i_gather_nw               (data_o_gather_nw[6][16]),
    .ready_o_gather_nw              (ready_i_gather_nw[6][16]),
    .valid_o_gather_nw              (valid_i_gather_nw[6][16]),
    .data_o_gather_nw               (data_i_gather_nw[6][16]),
    .ready_i_gather_nw              (ready_o_gather_nw[6][16]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[6][16]),
    .data_i_merge_nw                (data_o_merge_nw[6][16]),
    .ready_o_merge_nw               (ready_i_merge_nw[6][16]),
    .valid_o_merge_nw               (valid_i_merge_nw[6][16]),
    .data_o_merge_nw                (data_i_merge_nw[6][16]),
    .ready_i_merge_nw               (ready_o_merge_nw[6][16]),

    .valid_i_cast_pe                (cast_valid_i_6_16),
    .data_i_cast_pe                 (cast_data_i_6_16),
    .ready_o_cast_pe                (cast_ready_o_6_16),
    .valid_o_cast_pe                (cast_valid_o_6_16),
    .data_o_cast_pe                 (cast_data_o_6_16),
    .ready_i_cast_pe                (cast_ready_i_6_16),

    .valid_i_merge_pe               (merge_valid_i_6_16),
    .data_i_merge_pe                (merge_data_i_6_16),
    .ready_o_merge_pe               (merge_ready_o_6_16),
    .valid_o_merge_pe               (merge_valid_o_6_16),
    .data_o_merge_pe                (merge_data_o_6_16),
    .ready_i_merge_pe               (merge_ready_i_6_16),

    .valid_i_gather_pe              (gather_valid_i_6_16),
    .data_i_gather_pe               (gather_data_i_6_16),
    .ready_o_gather_pe              (gather_ready_o_6_16),
    .valid_o_gather_pe              (gather_valid_o_6_16),
    .data_o_gather_pe               (gather_data_o_6_16),
    .ready_i_gather_pe              (gather_ready_i_6_16),

    .credit_upd                     (credit_upd[6][16])
);


network_interface #(
    .cast_out                       (cast_out_6_17),
    .gather_out                     (gather_out_6_17),
    .cast_sid                       (cast_sid_6_17),
    .gather_sid                     (gather_sid_6_17)
)ni_6_17(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[6][17]),
    .data_i_cast_nw                 (data_o_cast_nw[6][17]),
    .ready_o_cast_nw                (ready_i_cast_nw[6][17]),
    .valid_o_cast_nw                (valid_i_cast_nw[6][17]),
    .data_o_cast_nw                 (data_i_cast_nw[6][17]),
    .ready_i_cast_nw                (ready_o_cast_nw[6][17]),

    .valid_i_gather_nw              (valid_o_gather_nw[6][17]),
    .data_i_gather_nw               (data_o_gather_nw[6][17]),
    .ready_o_gather_nw              (ready_i_gather_nw[6][17]),
    .valid_o_gather_nw              (valid_i_gather_nw[6][17]),
    .data_o_gather_nw               (data_i_gather_nw[6][17]),
    .ready_i_gather_nw              (ready_o_gather_nw[6][17]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[6][17]),
    .data_i_merge_nw                (data_o_merge_nw[6][17]),
    .ready_o_merge_nw               (ready_i_merge_nw[6][17]),
    .valid_o_merge_nw               (valid_i_merge_nw[6][17]),
    .data_o_merge_nw                (data_i_merge_nw[6][17]),
    .ready_i_merge_nw               (ready_o_merge_nw[6][17]),

    .valid_i_cast_pe                (cast_valid_i_6_17),
    .data_i_cast_pe                 (cast_data_i_6_17),
    .ready_o_cast_pe                (cast_ready_o_6_17),
    .valid_o_cast_pe                (cast_valid_o_6_17),
    .data_o_cast_pe                 (cast_data_o_6_17),
    .ready_i_cast_pe                (cast_ready_i_6_17),

    .valid_i_merge_pe               (merge_valid_i_6_17),
    .data_i_merge_pe                (merge_data_i_6_17),
    .ready_o_merge_pe               (merge_ready_o_6_17),
    .valid_o_merge_pe               (merge_valid_o_6_17),
    .data_o_merge_pe                (merge_data_o_6_17),
    .ready_i_merge_pe               (merge_ready_i_6_17),

    .valid_i_gather_pe              (gather_valid_i_6_17),
    .data_i_gather_pe               (gather_data_i_6_17),
    .ready_o_gather_pe              (gather_ready_o_6_17),
    .valid_o_gather_pe              (gather_valid_o_6_17),
    .data_o_gather_pe               (gather_data_o_6_17),
    .ready_i_gather_pe              (gather_ready_i_6_17),

    .credit_upd                     (credit_upd[6][17])
);


network_interface #(
    .cast_out                       (cast_out_6_18),
    .gather_out                     (gather_out_6_18),
    .cast_sid                       (cast_sid_6_18),
    .gather_sid                     (gather_sid_6_18)
)ni_6_18(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[6][18]),
    .data_i_cast_nw                 (data_o_cast_nw[6][18]),
    .ready_o_cast_nw                (ready_i_cast_nw[6][18]),
    .valid_o_cast_nw                (valid_i_cast_nw[6][18]),
    .data_o_cast_nw                 (data_i_cast_nw[6][18]),
    .ready_i_cast_nw                (ready_o_cast_nw[6][18]),

    .valid_i_gather_nw              (valid_o_gather_nw[6][18]),
    .data_i_gather_nw               (data_o_gather_nw[6][18]),
    .ready_o_gather_nw              (ready_i_gather_nw[6][18]),
    .valid_o_gather_nw              (valid_i_gather_nw[6][18]),
    .data_o_gather_nw               (data_i_gather_nw[6][18]),
    .ready_i_gather_nw              (ready_o_gather_nw[6][18]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[6][18]),
    .data_i_merge_nw                (data_o_merge_nw[6][18]),
    .ready_o_merge_nw               (ready_i_merge_nw[6][18]),
    .valid_o_merge_nw               (valid_i_merge_nw[6][18]),
    .data_o_merge_nw                (data_i_merge_nw[6][18]),
    .ready_i_merge_nw               (ready_o_merge_nw[6][18]),

    .valid_i_cast_pe                (cast_valid_i_6_18),
    .data_i_cast_pe                 (cast_data_i_6_18),
    .ready_o_cast_pe                (cast_ready_o_6_18),
    .valid_o_cast_pe                (cast_valid_o_6_18),
    .data_o_cast_pe                 (cast_data_o_6_18),
    .ready_i_cast_pe                (cast_ready_i_6_18),

    .valid_i_merge_pe               (merge_valid_i_6_18),
    .data_i_merge_pe                (merge_data_i_6_18),
    .ready_o_merge_pe               (merge_ready_o_6_18),
    .valid_o_merge_pe               (merge_valid_o_6_18),
    .data_o_merge_pe                (merge_data_o_6_18),
    .ready_i_merge_pe               (merge_ready_i_6_18),

    .valid_i_gather_pe              (gather_valid_i_6_18),
    .data_i_gather_pe               (gather_data_i_6_18),
    .ready_o_gather_pe              (gather_ready_o_6_18),
    .valid_o_gather_pe              (gather_valid_o_6_18),
    .data_o_gather_pe               (gather_data_o_6_18),
    .ready_i_gather_pe              (gather_ready_i_6_18),

    .credit_upd                     (credit_upd[6][18])
);


network_interface #(
    .cast_out                       (cast_out_6_19),
    .gather_out                     (gather_out_6_19),
    .cast_sid                       (cast_sid_6_19),
    .gather_sid                     (gather_sid_6_19)
)ni_6_19(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[6][19]),
    .data_i_cast_nw                 (data_o_cast_nw[6][19]),
    .ready_o_cast_nw                (ready_i_cast_nw[6][19]),
    .valid_o_cast_nw                (valid_i_cast_nw[6][19]),
    .data_o_cast_nw                 (data_i_cast_nw[6][19]),
    .ready_i_cast_nw                (ready_o_cast_nw[6][19]),

    .valid_i_gather_nw              (valid_o_gather_nw[6][19]),
    .data_i_gather_nw               (data_o_gather_nw[6][19]),
    .ready_o_gather_nw              (ready_i_gather_nw[6][19]),
    .valid_o_gather_nw              (valid_i_gather_nw[6][19]),
    .data_o_gather_nw               (data_i_gather_nw[6][19]),
    .ready_i_gather_nw              (ready_o_gather_nw[6][19]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[6][19]),
    .data_i_merge_nw                (data_o_merge_nw[6][19]),
    .ready_o_merge_nw               (ready_i_merge_nw[6][19]),
    .valid_o_merge_nw               (valid_i_merge_nw[6][19]),
    .data_o_merge_nw                (data_i_merge_nw[6][19]),
    .ready_i_merge_nw               (ready_o_merge_nw[6][19]),

    .valid_i_cast_pe                (cast_valid_i_6_19),
    .data_i_cast_pe                 (cast_data_i_6_19),
    .ready_o_cast_pe                (cast_ready_o_6_19),
    .valid_o_cast_pe                (cast_valid_o_6_19),
    .data_o_cast_pe                 (cast_data_o_6_19),
    .ready_i_cast_pe                (cast_ready_i_6_19),

    .valid_i_merge_pe               (merge_valid_i_6_19),
    .data_i_merge_pe                (merge_data_i_6_19),
    .ready_o_merge_pe               (merge_ready_o_6_19),
    .valid_o_merge_pe               (merge_valid_o_6_19),
    .data_o_merge_pe                (merge_data_o_6_19),
    .ready_i_merge_pe               (merge_ready_i_6_19),

    .valid_i_gather_pe              (gather_valid_i_6_19),
    .data_i_gather_pe               (gather_data_i_6_19),
    .ready_o_gather_pe              (gather_ready_o_6_19),
    .valid_o_gather_pe              (gather_valid_o_6_19),
    .data_o_gather_pe               (gather_data_o_6_19),
    .ready_i_gather_pe              (gather_ready_i_6_19),

    .credit_upd                     (credit_upd[6][19])
);


network_interface #(
    .cast_out                       (cast_out_6_20),
    .gather_out                     (gather_out_6_20),
    .cast_sid                       (cast_sid_6_20),
    .gather_sid                     (gather_sid_6_20)
)ni_6_20(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[6][20]),
    .data_i_cast_nw                 (data_o_cast_nw[6][20]),
    .ready_o_cast_nw                (ready_i_cast_nw[6][20]),
    .valid_o_cast_nw                (valid_i_cast_nw[6][20]),
    .data_o_cast_nw                 (data_i_cast_nw[6][20]),
    .ready_i_cast_nw                (ready_o_cast_nw[6][20]),

    .valid_i_gather_nw              (valid_o_gather_nw[6][20]),
    .data_i_gather_nw               (data_o_gather_nw[6][20]),
    .ready_o_gather_nw              (ready_i_gather_nw[6][20]),
    .valid_o_gather_nw              (valid_i_gather_nw[6][20]),
    .data_o_gather_nw               (data_i_gather_nw[6][20]),
    .ready_i_gather_nw              (ready_o_gather_nw[6][20]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[6][20]),
    .data_i_merge_nw                (data_o_merge_nw[6][20]),
    .ready_o_merge_nw               (ready_i_merge_nw[6][20]),
    .valid_o_merge_nw               (valid_i_merge_nw[6][20]),
    .data_o_merge_nw                (data_i_merge_nw[6][20]),
    .ready_i_merge_nw               (ready_o_merge_nw[6][20]),

    .valid_i_cast_pe                (cast_valid_i_6_20),
    .data_i_cast_pe                 (cast_data_i_6_20),
    .ready_o_cast_pe                (cast_ready_o_6_20),
    .valid_o_cast_pe                (cast_valid_o_6_20),
    .data_o_cast_pe                 (cast_data_o_6_20),
    .ready_i_cast_pe                (cast_ready_i_6_20),

    .valid_i_merge_pe               (merge_valid_i_6_20),
    .data_i_merge_pe                (merge_data_i_6_20),
    .ready_o_merge_pe               (merge_ready_o_6_20),
    .valid_o_merge_pe               (merge_valid_o_6_20),
    .data_o_merge_pe                (merge_data_o_6_20),
    .ready_i_merge_pe               (merge_ready_i_6_20),

    .valid_i_gather_pe              (gather_valid_i_6_20),
    .data_i_gather_pe               (gather_data_i_6_20),
    .ready_o_gather_pe              (gather_ready_o_6_20),
    .valid_o_gather_pe              (gather_valid_o_6_20),
    .data_o_gather_pe               (gather_data_o_6_20),
    .ready_i_gather_pe              (gather_ready_i_6_20),

    .credit_upd                     (credit_upd[6][20])
);


network_interface #(
    .cast_out                       (cast_out_6_21),
    .gather_out                     (gather_out_6_21),
    .cast_sid                       (cast_sid_6_21),
    .gather_sid                     (gather_sid_6_21)
)ni_6_21(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[6][21]),
    .data_i_cast_nw                 (data_o_cast_nw[6][21]),
    .ready_o_cast_nw                (ready_i_cast_nw[6][21]),
    .valid_o_cast_nw                (valid_i_cast_nw[6][21]),
    .data_o_cast_nw                 (data_i_cast_nw[6][21]),
    .ready_i_cast_nw                (ready_o_cast_nw[6][21]),

    .valid_i_gather_nw              (valid_o_gather_nw[6][21]),
    .data_i_gather_nw               (data_o_gather_nw[6][21]),
    .ready_o_gather_nw              (ready_i_gather_nw[6][21]),
    .valid_o_gather_nw              (valid_i_gather_nw[6][21]),
    .data_o_gather_nw               (data_i_gather_nw[6][21]),
    .ready_i_gather_nw              (ready_o_gather_nw[6][21]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[6][21]),
    .data_i_merge_nw                (data_o_merge_nw[6][21]),
    .ready_o_merge_nw               (ready_i_merge_nw[6][21]),
    .valid_o_merge_nw               (valid_i_merge_nw[6][21]),
    .data_o_merge_nw                (data_i_merge_nw[6][21]),
    .ready_i_merge_nw               (ready_o_merge_nw[6][21]),

    .valid_i_cast_pe                (cast_valid_i_6_21),
    .data_i_cast_pe                 (cast_data_i_6_21),
    .ready_o_cast_pe                (cast_ready_o_6_21),
    .valid_o_cast_pe                (cast_valid_o_6_21),
    .data_o_cast_pe                 (cast_data_o_6_21),
    .ready_i_cast_pe                (cast_ready_i_6_21),

    .valid_i_merge_pe               (merge_valid_i_6_21),
    .data_i_merge_pe                (merge_data_i_6_21),
    .ready_o_merge_pe               (merge_ready_o_6_21),
    .valid_o_merge_pe               (merge_valid_o_6_21),
    .data_o_merge_pe                (merge_data_o_6_21),
    .ready_i_merge_pe               (merge_ready_i_6_21),

    .valid_i_gather_pe              (gather_valid_i_6_21),
    .data_i_gather_pe               (gather_data_i_6_21),
    .ready_o_gather_pe              (gather_ready_o_6_21),
    .valid_o_gather_pe              (gather_valid_o_6_21),
    .data_o_gather_pe               (gather_data_o_6_21),
    .ready_i_gather_pe              (gather_ready_i_6_21),

    .credit_upd                     (credit_upd[6][21])
);


network_interface #(
    .cast_out                       (cast_out_6_22),
    .gather_out                     (gather_out_6_22),
    .cast_sid                       (cast_sid_6_22),
    .gather_sid                     (gather_sid_6_22)
)ni_6_22(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[6][22]),
    .data_i_cast_nw                 (data_o_cast_nw[6][22]),
    .ready_o_cast_nw                (ready_i_cast_nw[6][22]),
    .valid_o_cast_nw                (valid_i_cast_nw[6][22]),
    .data_o_cast_nw                 (data_i_cast_nw[6][22]),
    .ready_i_cast_nw                (ready_o_cast_nw[6][22]),

    .valid_i_gather_nw              (valid_o_gather_nw[6][22]),
    .data_i_gather_nw               (data_o_gather_nw[6][22]),
    .ready_o_gather_nw              (ready_i_gather_nw[6][22]),
    .valid_o_gather_nw              (valid_i_gather_nw[6][22]),
    .data_o_gather_nw               (data_i_gather_nw[6][22]),
    .ready_i_gather_nw              (ready_o_gather_nw[6][22]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[6][22]),
    .data_i_merge_nw                (data_o_merge_nw[6][22]),
    .ready_o_merge_nw               (ready_i_merge_nw[6][22]),
    .valid_o_merge_nw               (valid_i_merge_nw[6][22]),
    .data_o_merge_nw                (data_i_merge_nw[6][22]),
    .ready_i_merge_nw               (ready_o_merge_nw[6][22]),

    .valid_i_cast_pe                (cast_valid_i_6_22),
    .data_i_cast_pe                 (cast_data_i_6_22),
    .ready_o_cast_pe                (cast_ready_o_6_22),
    .valid_o_cast_pe                (cast_valid_o_6_22),
    .data_o_cast_pe                 (cast_data_o_6_22),
    .ready_i_cast_pe                (cast_ready_i_6_22),

    .valid_i_merge_pe               (merge_valid_i_6_22),
    .data_i_merge_pe                (merge_data_i_6_22),
    .ready_o_merge_pe               (merge_ready_o_6_22),
    .valid_o_merge_pe               (merge_valid_o_6_22),
    .data_o_merge_pe                (merge_data_o_6_22),
    .ready_i_merge_pe               (merge_ready_i_6_22),

    .valid_i_gather_pe              (gather_valid_i_6_22),
    .data_i_gather_pe               (gather_data_i_6_22),
    .ready_o_gather_pe              (gather_ready_o_6_22),
    .valid_o_gather_pe              (gather_valid_o_6_22),
    .data_o_gather_pe               (gather_data_o_6_22),
    .ready_i_gather_pe              (gather_ready_i_6_22),

    .credit_upd                     (credit_upd[6][22])
);


network_interface #(
    .cast_out                       (cast_out_6_23),
    .gather_out                     (gather_out_6_23),
    .cast_sid                       (cast_sid_6_23),
    .gather_sid                     (gather_sid_6_23)
)ni_6_23(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[6][23]),
    .data_i_cast_nw                 (data_o_cast_nw[6][23]),
    .ready_o_cast_nw                (ready_i_cast_nw[6][23]),
    .valid_o_cast_nw                (valid_i_cast_nw[6][23]),
    .data_o_cast_nw                 (data_i_cast_nw[6][23]),
    .ready_i_cast_nw                (ready_o_cast_nw[6][23]),

    .valid_i_gather_nw              (valid_o_gather_nw[6][23]),
    .data_i_gather_nw               (data_o_gather_nw[6][23]),
    .ready_o_gather_nw              (ready_i_gather_nw[6][23]),
    .valid_o_gather_nw              (valid_i_gather_nw[6][23]),
    .data_o_gather_nw               (data_i_gather_nw[6][23]),
    .ready_i_gather_nw              (ready_o_gather_nw[6][23]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[6][23]),
    .data_i_merge_nw                (data_o_merge_nw[6][23]),
    .ready_o_merge_nw               (ready_i_merge_nw[6][23]),
    .valid_o_merge_nw               (valid_i_merge_nw[6][23]),
    .data_o_merge_nw                (data_i_merge_nw[6][23]),
    .ready_i_merge_nw               (ready_o_merge_nw[6][23]),

    .valid_i_cast_pe                (cast_valid_i_6_23),
    .data_i_cast_pe                 (cast_data_i_6_23),
    .ready_o_cast_pe                (cast_ready_o_6_23),
    .valid_o_cast_pe                (cast_valid_o_6_23),
    .data_o_cast_pe                 (cast_data_o_6_23),
    .ready_i_cast_pe                (cast_ready_i_6_23),

    .valid_i_merge_pe               (merge_valid_i_6_23),
    .data_i_merge_pe                (merge_data_i_6_23),
    .ready_o_merge_pe               (merge_ready_o_6_23),
    .valid_o_merge_pe               (merge_valid_o_6_23),
    .data_o_merge_pe                (merge_data_o_6_23),
    .ready_i_merge_pe               (merge_ready_i_6_23),

    .valid_i_gather_pe              (gather_valid_i_6_23),
    .data_i_gather_pe               (gather_data_i_6_23),
    .ready_o_gather_pe              (gather_ready_o_6_23),
    .valid_o_gather_pe              (gather_valid_o_6_23),
    .data_o_gather_pe               (gather_data_o_6_23),
    .ready_i_gather_pe              (gather_ready_i_6_23),

    .credit_upd                     (credit_upd[6][23])
);


network_interface #(
    .cast_out                       (cast_out_6_24),
    .gather_out                     (gather_out_6_24),
    .cast_sid                       (cast_sid_6_24),
    .gather_sid                     (gather_sid_6_24)
)ni_6_24(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[6][24]),
    .data_i_cast_nw                 (data_o_cast_nw[6][24]),
    .ready_o_cast_nw                (ready_i_cast_nw[6][24]),
    .valid_o_cast_nw                (valid_i_cast_nw[6][24]),
    .data_o_cast_nw                 (data_i_cast_nw[6][24]),
    .ready_i_cast_nw                (ready_o_cast_nw[6][24]),

    .valid_i_gather_nw              (valid_o_gather_nw[6][24]),
    .data_i_gather_nw               (data_o_gather_nw[6][24]),
    .ready_o_gather_nw              (ready_i_gather_nw[6][24]),
    .valid_o_gather_nw              (valid_i_gather_nw[6][24]),
    .data_o_gather_nw               (data_i_gather_nw[6][24]),
    .ready_i_gather_nw              (ready_o_gather_nw[6][24]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[6][24]),
    .data_i_merge_nw                (data_o_merge_nw[6][24]),
    .ready_o_merge_nw               (ready_i_merge_nw[6][24]),
    .valid_o_merge_nw               (valid_i_merge_nw[6][24]),
    .data_o_merge_nw                (data_i_merge_nw[6][24]),
    .ready_i_merge_nw               (ready_o_merge_nw[6][24]),

    .valid_i_cast_pe                (cast_valid_i_6_24),
    .data_i_cast_pe                 (cast_data_i_6_24),
    .ready_o_cast_pe                (cast_ready_o_6_24),
    .valid_o_cast_pe                (cast_valid_o_6_24),
    .data_o_cast_pe                 (cast_data_o_6_24),
    .ready_i_cast_pe                (cast_ready_i_6_24),

    .valid_i_merge_pe               (merge_valid_i_6_24),
    .data_i_merge_pe                (merge_data_i_6_24),
    .ready_o_merge_pe               (merge_ready_o_6_24),
    .valid_o_merge_pe               (merge_valid_o_6_24),
    .data_o_merge_pe                (merge_data_o_6_24),
    .ready_i_merge_pe               (merge_ready_i_6_24),

    .valid_i_gather_pe              (gather_valid_i_6_24),
    .data_i_gather_pe               (gather_data_i_6_24),
    .ready_o_gather_pe              (gather_ready_o_6_24),
    .valid_o_gather_pe              (gather_valid_o_6_24),
    .data_o_gather_pe               (gather_data_o_6_24),
    .ready_i_gather_pe              (gather_ready_i_6_24),

    .credit_upd                     (credit_upd[6][24])
);


network_interface #(
    .cast_out                       (cast_out_7_0),
    .gather_out                     (gather_out_7_0),
    .cast_sid                       (cast_sid_7_0),
    .gather_sid                     (gather_sid_7_0)
)ni_7_0(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[7][0]),
    .data_i_cast_nw                 (data_o_cast_nw[7][0]),
    .ready_o_cast_nw                (ready_i_cast_nw[7][0]),
    .valid_o_cast_nw                (valid_i_cast_nw[7][0]),
    .data_o_cast_nw                 (data_i_cast_nw[7][0]),
    .ready_i_cast_nw                (ready_o_cast_nw[7][0]),

    .valid_i_gather_nw              (valid_o_gather_nw[7][0]),
    .data_i_gather_nw               (data_o_gather_nw[7][0]),
    .ready_o_gather_nw              (ready_i_gather_nw[7][0]),
    .valid_o_gather_nw              (valid_i_gather_nw[7][0]),
    .data_o_gather_nw               (data_i_gather_nw[7][0]),
    .ready_i_gather_nw              (ready_o_gather_nw[7][0]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[7][0]),
    .data_i_merge_nw                (data_o_merge_nw[7][0]),
    .ready_o_merge_nw               (ready_i_merge_nw[7][0]),
    .valid_o_merge_nw               (valid_i_merge_nw[7][0]),
    .data_o_merge_nw                (data_i_merge_nw[7][0]),
    .ready_i_merge_nw               (ready_o_merge_nw[7][0]),

    .valid_i_cast_pe                (cast_valid_i_7_0),
    .data_i_cast_pe                 (cast_data_i_7_0),
    .ready_o_cast_pe                (cast_ready_o_7_0),
    .valid_o_cast_pe                (cast_valid_o_7_0),
    .data_o_cast_pe                 (cast_data_o_7_0),
    .ready_i_cast_pe                (cast_ready_i_7_0),

    .valid_i_merge_pe               (merge_valid_i_7_0),
    .data_i_merge_pe                (merge_data_i_7_0),
    .ready_o_merge_pe               (merge_ready_o_7_0),
    .valid_o_merge_pe               (merge_valid_o_7_0),
    .data_o_merge_pe                (merge_data_o_7_0),
    .ready_i_merge_pe               (merge_ready_i_7_0),

    .valid_i_gather_pe              (gather_valid_i_7_0),
    .data_i_gather_pe               (gather_data_i_7_0),
    .ready_o_gather_pe              (gather_ready_o_7_0),
    .valid_o_gather_pe              (gather_valid_o_7_0),
    .data_o_gather_pe               (gather_data_o_7_0),
    .ready_i_gather_pe              (gather_ready_i_7_0),

    .credit_upd                     (credit_upd[7][0])
);


network_interface #(
    .cast_out                       (cast_out_7_1),
    .gather_out                     (gather_out_7_1),
    .cast_sid                       (cast_sid_7_1),
    .gather_sid                     (gather_sid_7_1)
)ni_7_1(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[7][1]),
    .data_i_cast_nw                 (data_o_cast_nw[7][1]),
    .ready_o_cast_nw                (ready_i_cast_nw[7][1]),
    .valid_o_cast_nw                (valid_i_cast_nw[7][1]),
    .data_o_cast_nw                 (data_i_cast_nw[7][1]),
    .ready_i_cast_nw                (ready_o_cast_nw[7][1]),

    .valid_i_gather_nw              (valid_o_gather_nw[7][1]),
    .data_i_gather_nw               (data_o_gather_nw[7][1]),
    .ready_o_gather_nw              (ready_i_gather_nw[7][1]),
    .valid_o_gather_nw              (valid_i_gather_nw[7][1]),
    .data_o_gather_nw               (data_i_gather_nw[7][1]),
    .ready_i_gather_nw              (ready_o_gather_nw[7][1]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[7][1]),
    .data_i_merge_nw                (data_o_merge_nw[7][1]),
    .ready_o_merge_nw               (ready_i_merge_nw[7][1]),
    .valid_o_merge_nw               (valid_i_merge_nw[7][1]),
    .data_o_merge_nw                (data_i_merge_nw[7][1]),
    .ready_i_merge_nw               (ready_o_merge_nw[7][1]),

    .valid_i_cast_pe                (cast_valid_i_7_1),
    .data_i_cast_pe                 (cast_data_i_7_1),
    .ready_o_cast_pe                (cast_ready_o_7_1),
    .valid_o_cast_pe                (cast_valid_o_7_1),
    .data_o_cast_pe                 (cast_data_o_7_1),
    .ready_i_cast_pe                (cast_ready_i_7_1),

    .valid_i_merge_pe               (merge_valid_i_7_1),
    .data_i_merge_pe                (merge_data_i_7_1),
    .ready_o_merge_pe               (merge_ready_o_7_1),
    .valid_o_merge_pe               (merge_valid_o_7_1),
    .data_o_merge_pe                (merge_data_o_7_1),
    .ready_i_merge_pe               (merge_ready_i_7_1),

    .valid_i_gather_pe              (gather_valid_i_7_1),
    .data_i_gather_pe               (gather_data_i_7_1),
    .ready_o_gather_pe              (gather_ready_o_7_1),
    .valid_o_gather_pe              (gather_valid_o_7_1),
    .data_o_gather_pe               (gather_data_o_7_1),
    .ready_i_gather_pe              (gather_ready_i_7_1),

    .credit_upd                     (credit_upd[7][1])
);


network_interface #(
    .cast_out                       (cast_out_7_2),
    .gather_out                     (gather_out_7_2),
    .cast_sid                       (cast_sid_7_2),
    .gather_sid                     (gather_sid_7_2)
)ni_7_2(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[7][2]),
    .data_i_cast_nw                 (data_o_cast_nw[7][2]),
    .ready_o_cast_nw                (ready_i_cast_nw[7][2]),
    .valid_o_cast_nw                (valid_i_cast_nw[7][2]),
    .data_o_cast_nw                 (data_i_cast_nw[7][2]),
    .ready_i_cast_nw                (ready_o_cast_nw[7][2]),

    .valid_i_gather_nw              (valid_o_gather_nw[7][2]),
    .data_i_gather_nw               (data_o_gather_nw[7][2]),
    .ready_o_gather_nw              (ready_i_gather_nw[7][2]),
    .valid_o_gather_nw              (valid_i_gather_nw[7][2]),
    .data_o_gather_nw               (data_i_gather_nw[7][2]),
    .ready_i_gather_nw              (ready_o_gather_nw[7][2]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[7][2]),
    .data_i_merge_nw                (data_o_merge_nw[7][2]),
    .ready_o_merge_nw               (ready_i_merge_nw[7][2]),
    .valid_o_merge_nw               (valid_i_merge_nw[7][2]),
    .data_o_merge_nw                (data_i_merge_nw[7][2]),
    .ready_i_merge_nw               (ready_o_merge_nw[7][2]),

    .valid_i_cast_pe                (cast_valid_i_7_2),
    .data_i_cast_pe                 (cast_data_i_7_2),
    .ready_o_cast_pe                (cast_ready_o_7_2),
    .valid_o_cast_pe                (cast_valid_o_7_2),
    .data_o_cast_pe                 (cast_data_o_7_2),
    .ready_i_cast_pe                (cast_ready_i_7_2),

    .valid_i_merge_pe               (merge_valid_i_7_2),
    .data_i_merge_pe                (merge_data_i_7_2),
    .ready_o_merge_pe               (merge_ready_o_7_2),
    .valid_o_merge_pe               (merge_valid_o_7_2),
    .data_o_merge_pe                (merge_data_o_7_2),
    .ready_i_merge_pe               (merge_ready_i_7_2),

    .valid_i_gather_pe              (gather_valid_i_7_2),
    .data_i_gather_pe               (gather_data_i_7_2),
    .ready_o_gather_pe              (gather_ready_o_7_2),
    .valid_o_gather_pe              (gather_valid_o_7_2),
    .data_o_gather_pe               (gather_data_o_7_2),
    .ready_i_gather_pe              (gather_ready_i_7_2),

    .credit_upd                     (credit_upd[7][2])
);


network_interface #(
    .cast_out                       (cast_out_7_3),
    .gather_out                     (gather_out_7_3),
    .cast_sid                       (cast_sid_7_3),
    .gather_sid                     (gather_sid_7_3)
)ni_7_3(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[7][3]),
    .data_i_cast_nw                 (data_o_cast_nw[7][3]),
    .ready_o_cast_nw                (ready_i_cast_nw[7][3]),
    .valid_o_cast_nw                (valid_i_cast_nw[7][3]),
    .data_o_cast_nw                 (data_i_cast_nw[7][3]),
    .ready_i_cast_nw                (ready_o_cast_nw[7][3]),

    .valid_i_gather_nw              (valid_o_gather_nw[7][3]),
    .data_i_gather_nw               (data_o_gather_nw[7][3]),
    .ready_o_gather_nw              (ready_i_gather_nw[7][3]),
    .valid_o_gather_nw              (valid_i_gather_nw[7][3]),
    .data_o_gather_nw               (data_i_gather_nw[7][3]),
    .ready_i_gather_nw              (ready_o_gather_nw[7][3]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[7][3]),
    .data_i_merge_nw                (data_o_merge_nw[7][3]),
    .ready_o_merge_nw               (ready_i_merge_nw[7][3]),
    .valid_o_merge_nw               (valid_i_merge_nw[7][3]),
    .data_o_merge_nw                (data_i_merge_nw[7][3]),
    .ready_i_merge_nw               (ready_o_merge_nw[7][3]),

    .valid_i_cast_pe                (cast_valid_i_7_3),
    .data_i_cast_pe                 (cast_data_i_7_3),
    .ready_o_cast_pe                (cast_ready_o_7_3),
    .valid_o_cast_pe                (cast_valid_o_7_3),
    .data_o_cast_pe                 (cast_data_o_7_3),
    .ready_i_cast_pe                (cast_ready_i_7_3),

    .valid_i_merge_pe               (merge_valid_i_7_3),
    .data_i_merge_pe                (merge_data_i_7_3),
    .ready_o_merge_pe               (merge_ready_o_7_3),
    .valid_o_merge_pe               (merge_valid_o_7_3),
    .data_o_merge_pe                (merge_data_o_7_3),
    .ready_i_merge_pe               (merge_ready_i_7_3),

    .valid_i_gather_pe              (gather_valid_i_7_3),
    .data_i_gather_pe               (gather_data_i_7_3),
    .ready_o_gather_pe              (gather_ready_o_7_3),
    .valid_o_gather_pe              (gather_valid_o_7_3),
    .data_o_gather_pe               (gather_data_o_7_3),
    .ready_i_gather_pe              (gather_ready_i_7_3),

    .credit_upd                     (credit_upd[7][3])
);


network_interface #(
    .cast_out                       (cast_out_7_4),
    .gather_out                     (gather_out_7_4),
    .cast_sid                       (cast_sid_7_4),
    .gather_sid                     (gather_sid_7_4)
)ni_7_4(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[7][4]),
    .data_i_cast_nw                 (data_o_cast_nw[7][4]),
    .ready_o_cast_nw                (ready_i_cast_nw[7][4]),
    .valid_o_cast_nw                (valid_i_cast_nw[7][4]),
    .data_o_cast_nw                 (data_i_cast_nw[7][4]),
    .ready_i_cast_nw                (ready_o_cast_nw[7][4]),

    .valid_i_gather_nw              (valid_o_gather_nw[7][4]),
    .data_i_gather_nw               (data_o_gather_nw[7][4]),
    .ready_o_gather_nw              (ready_i_gather_nw[7][4]),
    .valid_o_gather_nw              (valid_i_gather_nw[7][4]),
    .data_o_gather_nw               (data_i_gather_nw[7][4]),
    .ready_i_gather_nw              (ready_o_gather_nw[7][4]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[7][4]),
    .data_i_merge_nw                (data_o_merge_nw[7][4]),
    .ready_o_merge_nw               (ready_i_merge_nw[7][4]),
    .valid_o_merge_nw               (valid_i_merge_nw[7][4]),
    .data_o_merge_nw                (data_i_merge_nw[7][4]),
    .ready_i_merge_nw               (ready_o_merge_nw[7][4]),

    .valid_i_cast_pe                (cast_valid_i_7_4),
    .data_i_cast_pe                 (cast_data_i_7_4),
    .ready_o_cast_pe                (cast_ready_o_7_4),
    .valid_o_cast_pe                (cast_valid_o_7_4),
    .data_o_cast_pe                 (cast_data_o_7_4),
    .ready_i_cast_pe                (cast_ready_i_7_4),

    .valid_i_merge_pe               (merge_valid_i_7_4),
    .data_i_merge_pe                (merge_data_i_7_4),
    .ready_o_merge_pe               (merge_ready_o_7_4),
    .valid_o_merge_pe               (merge_valid_o_7_4),
    .data_o_merge_pe                (merge_data_o_7_4),
    .ready_i_merge_pe               (merge_ready_i_7_4),

    .valid_i_gather_pe              (gather_valid_i_7_4),
    .data_i_gather_pe               (gather_data_i_7_4),
    .ready_o_gather_pe              (gather_ready_o_7_4),
    .valid_o_gather_pe              (gather_valid_o_7_4),
    .data_o_gather_pe               (gather_data_o_7_4),
    .ready_i_gather_pe              (gather_ready_i_7_4),

    .credit_upd                     (credit_upd[7][4])
);


network_interface #(
    .cast_out                       (cast_out_7_5),
    .gather_out                     (gather_out_7_5),
    .cast_sid                       (cast_sid_7_5),
    .gather_sid                     (gather_sid_7_5)
)ni_7_5(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[7][5]),
    .data_i_cast_nw                 (data_o_cast_nw[7][5]),
    .ready_o_cast_nw                (ready_i_cast_nw[7][5]),
    .valid_o_cast_nw                (valid_i_cast_nw[7][5]),
    .data_o_cast_nw                 (data_i_cast_nw[7][5]),
    .ready_i_cast_nw                (ready_o_cast_nw[7][5]),

    .valid_i_gather_nw              (valid_o_gather_nw[7][5]),
    .data_i_gather_nw               (data_o_gather_nw[7][5]),
    .ready_o_gather_nw              (ready_i_gather_nw[7][5]),
    .valid_o_gather_nw              (valid_i_gather_nw[7][5]),
    .data_o_gather_nw               (data_i_gather_nw[7][5]),
    .ready_i_gather_nw              (ready_o_gather_nw[7][5]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[7][5]),
    .data_i_merge_nw                (data_o_merge_nw[7][5]),
    .ready_o_merge_nw               (ready_i_merge_nw[7][5]),
    .valid_o_merge_nw               (valid_i_merge_nw[7][5]),
    .data_o_merge_nw                (data_i_merge_nw[7][5]),
    .ready_i_merge_nw               (ready_o_merge_nw[7][5]),

    .valid_i_cast_pe                (cast_valid_i_7_5),
    .data_i_cast_pe                 (cast_data_i_7_5),
    .ready_o_cast_pe                (cast_ready_o_7_5),
    .valid_o_cast_pe                (cast_valid_o_7_5),
    .data_o_cast_pe                 (cast_data_o_7_5),
    .ready_i_cast_pe                (cast_ready_i_7_5),

    .valid_i_merge_pe               (merge_valid_i_7_5),
    .data_i_merge_pe                (merge_data_i_7_5),
    .ready_o_merge_pe               (merge_ready_o_7_5),
    .valid_o_merge_pe               (merge_valid_o_7_5),
    .data_o_merge_pe                (merge_data_o_7_5),
    .ready_i_merge_pe               (merge_ready_i_7_5),

    .valid_i_gather_pe              (gather_valid_i_7_5),
    .data_i_gather_pe               (gather_data_i_7_5),
    .ready_o_gather_pe              (gather_ready_o_7_5),
    .valid_o_gather_pe              (gather_valid_o_7_5),
    .data_o_gather_pe               (gather_data_o_7_5),
    .ready_i_gather_pe              (gather_ready_i_7_5),

    .credit_upd                     (credit_upd[7][5])
);


network_interface #(
    .cast_out                       (cast_out_7_6),
    .gather_out                     (gather_out_7_6),
    .cast_sid                       (cast_sid_7_6),
    .gather_sid                     (gather_sid_7_6)
)ni_7_6(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[7][6]),
    .data_i_cast_nw                 (data_o_cast_nw[7][6]),
    .ready_o_cast_nw                (ready_i_cast_nw[7][6]),
    .valid_o_cast_nw                (valid_i_cast_nw[7][6]),
    .data_o_cast_nw                 (data_i_cast_nw[7][6]),
    .ready_i_cast_nw                (ready_o_cast_nw[7][6]),

    .valid_i_gather_nw              (valid_o_gather_nw[7][6]),
    .data_i_gather_nw               (data_o_gather_nw[7][6]),
    .ready_o_gather_nw              (ready_i_gather_nw[7][6]),
    .valid_o_gather_nw              (valid_i_gather_nw[7][6]),
    .data_o_gather_nw               (data_i_gather_nw[7][6]),
    .ready_i_gather_nw              (ready_o_gather_nw[7][6]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[7][6]),
    .data_i_merge_nw                (data_o_merge_nw[7][6]),
    .ready_o_merge_nw               (ready_i_merge_nw[7][6]),
    .valid_o_merge_nw               (valid_i_merge_nw[7][6]),
    .data_o_merge_nw                (data_i_merge_nw[7][6]),
    .ready_i_merge_nw               (ready_o_merge_nw[7][6]),

    .valid_i_cast_pe                (cast_valid_i_7_6),
    .data_i_cast_pe                 (cast_data_i_7_6),
    .ready_o_cast_pe                (cast_ready_o_7_6),
    .valid_o_cast_pe                (cast_valid_o_7_6),
    .data_o_cast_pe                 (cast_data_o_7_6),
    .ready_i_cast_pe                (cast_ready_i_7_6),

    .valid_i_merge_pe               (merge_valid_i_7_6),
    .data_i_merge_pe                (merge_data_i_7_6),
    .ready_o_merge_pe               (merge_ready_o_7_6),
    .valid_o_merge_pe               (merge_valid_o_7_6),
    .data_o_merge_pe                (merge_data_o_7_6),
    .ready_i_merge_pe               (merge_ready_i_7_6),

    .valid_i_gather_pe              (gather_valid_i_7_6),
    .data_i_gather_pe               (gather_data_i_7_6),
    .ready_o_gather_pe              (gather_ready_o_7_6),
    .valid_o_gather_pe              (gather_valid_o_7_6),
    .data_o_gather_pe               (gather_data_o_7_6),
    .ready_i_gather_pe              (gather_ready_i_7_6),

    .credit_upd                     (credit_upd[7][6])
);


network_interface #(
    .cast_out                       (cast_out_7_7),
    .gather_out                     (gather_out_7_7),
    .cast_sid                       (cast_sid_7_7),
    .gather_sid                     (gather_sid_7_7)
)ni_7_7(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[7][7]),
    .data_i_cast_nw                 (data_o_cast_nw[7][7]),
    .ready_o_cast_nw                (ready_i_cast_nw[7][7]),
    .valid_o_cast_nw                (valid_i_cast_nw[7][7]),
    .data_o_cast_nw                 (data_i_cast_nw[7][7]),
    .ready_i_cast_nw                (ready_o_cast_nw[7][7]),

    .valid_i_gather_nw              (valid_o_gather_nw[7][7]),
    .data_i_gather_nw               (data_o_gather_nw[7][7]),
    .ready_o_gather_nw              (ready_i_gather_nw[7][7]),
    .valid_o_gather_nw              (valid_i_gather_nw[7][7]),
    .data_o_gather_nw               (data_i_gather_nw[7][7]),
    .ready_i_gather_nw              (ready_o_gather_nw[7][7]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[7][7]),
    .data_i_merge_nw                (data_o_merge_nw[7][7]),
    .ready_o_merge_nw               (ready_i_merge_nw[7][7]),
    .valid_o_merge_nw               (valid_i_merge_nw[7][7]),
    .data_o_merge_nw                (data_i_merge_nw[7][7]),
    .ready_i_merge_nw               (ready_o_merge_nw[7][7]),

    .valid_i_cast_pe                (cast_valid_i_7_7),
    .data_i_cast_pe                 (cast_data_i_7_7),
    .ready_o_cast_pe                (cast_ready_o_7_7),
    .valid_o_cast_pe                (cast_valid_o_7_7),
    .data_o_cast_pe                 (cast_data_o_7_7),
    .ready_i_cast_pe                (cast_ready_i_7_7),

    .valid_i_merge_pe               (merge_valid_i_7_7),
    .data_i_merge_pe                (merge_data_i_7_7),
    .ready_o_merge_pe               (merge_ready_o_7_7),
    .valid_o_merge_pe               (merge_valid_o_7_7),
    .data_o_merge_pe                (merge_data_o_7_7),
    .ready_i_merge_pe               (merge_ready_i_7_7),

    .valid_i_gather_pe              (gather_valid_i_7_7),
    .data_i_gather_pe               (gather_data_i_7_7),
    .ready_o_gather_pe              (gather_ready_o_7_7),
    .valid_o_gather_pe              (gather_valid_o_7_7),
    .data_o_gather_pe               (gather_data_o_7_7),
    .ready_i_gather_pe              (gather_ready_i_7_7),

    .credit_upd                     (credit_upd[7][7])
);


network_interface #(
    .cast_out                       (cast_out_7_8),
    .gather_out                     (gather_out_7_8),
    .cast_sid                       (cast_sid_7_8),
    .gather_sid                     (gather_sid_7_8)
)ni_7_8(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[7][8]),
    .data_i_cast_nw                 (data_o_cast_nw[7][8]),
    .ready_o_cast_nw                (ready_i_cast_nw[7][8]),
    .valid_o_cast_nw                (valid_i_cast_nw[7][8]),
    .data_o_cast_nw                 (data_i_cast_nw[7][8]),
    .ready_i_cast_nw                (ready_o_cast_nw[7][8]),

    .valid_i_gather_nw              (valid_o_gather_nw[7][8]),
    .data_i_gather_nw               (data_o_gather_nw[7][8]),
    .ready_o_gather_nw              (ready_i_gather_nw[7][8]),
    .valid_o_gather_nw              (valid_i_gather_nw[7][8]),
    .data_o_gather_nw               (data_i_gather_nw[7][8]),
    .ready_i_gather_nw              (ready_o_gather_nw[7][8]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[7][8]),
    .data_i_merge_nw                (data_o_merge_nw[7][8]),
    .ready_o_merge_nw               (ready_i_merge_nw[7][8]),
    .valid_o_merge_nw               (valid_i_merge_nw[7][8]),
    .data_o_merge_nw                (data_i_merge_nw[7][8]),
    .ready_i_merge_nw               (ready_o_merge_nw[7][8]),

    .valid_i_cast_pe                (cast_valid_i_7_8),
    .data_i_cast_pe                 (cast_data_i_7_8),
    .ready_o_cast_pe                (cast_ready_o_7_8),
    .valid_o_cast_pe                (cast_valid_o_7_8),
    .data_o_cast_pe                 (cast_data_o_7_8),
    .ready_i_cast_pe                (cast_ready_i_7_8),

    .valid_i_merge_pe               (merge_valid_i_7_8),
    .data_i_merge_pe                (merge_data_i_7_8),
    .ready_o_merge_pe               (merge_ready_o_7_8),
    .valid_o_merge_pe               (merge_valid_o_7_8),
    .data_o_merge_pe                (merge_data_o_7_8),
    .ready_i_merge_pe               (merge_ready_i_7_8),

    .valid_i_gather_pe              (gather_valid_i_7_8),
    .data_i_gather_pe               (gather_data_i_7_8),
    .ready_o_gather_pe              (gather_ready_o_7_8),
    .valid_o_gather_pe              (gather_valid_o_7_8),
    .data_o_gather_pe               (gather_data_o_7_8),
    .ready_i_gather_pe              (gather_ready_i_7_8),

    .credit_upd                     (credit_upd[7][8])
);


network_interface #(
    .cast_out                       (cast_out_7_9),
    .gather_out                     (gather_out_7_9),
    .cast_sid                       (cast_sid_7_9),
    .gather_sid                     (gather_sid_7_9)
)ni_7_9(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[7][9]),
    .data_i_cast_nw                 (data_o_cast_nw[7][9]),
    .ready_o_cast_nw                (ready_i_cast_nw[7][9]),
    .valid_o_cast_nw                (valid_i_cast_nw[7][9]),
    .data_o_cast_nw                 (data_i_cast_nw[7][9]),
    .ready_i_cast_nw                (ready_o_cast_nw[7][9]),

    .valid_i_gather_nw              (valid_o_gather_nw[7][9]),
    .data_i_gather_nw               (data_o_gather_nw[7][9]),
    .ready_o_gather_nw              (ready_i_gather_nw[7][9]),
    .valid_o_gather_nw              (valid_i_gather_nw[7][9]),
    .data_o_gather_nw               (data_i_gather_nw[7][9]),
    .ready_i_gather_nw              (ready_o_gather_nw[7][9]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[7][9]),
    .data_i_merge_nw                (data_o_merge_nw[7][9]),
    .ready_o_merge_nw               (ready_i_merge_nw[7][9]),
    .valid_o_merge_nw               (valid_i_merge_nw[7][9]),
    .data_o_merge_nw                (data_i_merge_nw[7][9]),
    .ready_i_merge_nw               (ready_o_merge_nw[7][9]),

    .valid_i_cast_pe                (cast_valid_i_7_9),
    .data_i_cast_pe                 (cast_data_i_7_9),
    .ready_o_cast_pe                (cast_ready_o_7_9),
    .valid_o_cast_pe                (cast_valid_o_7_9),
    .data_o_cast_pe                 (cast_data_o_7_9),
    .ready_i_cast_pe                (cast_ready_i_7_9),

    .valid_i_merge_pe               (merge_valid_i_7_9),
    .data_i_merge_pe                (merge_data_i_7_9),
    .ready_o_merge_pe               (merge_ready_o_7_9),
    .valid_o_merge_pe               (merge_valid_o_7_9),
    .data_o_merge_pe                (merge_data_o_7_9),
    .ready_i_merge_pe               (merge_ready_i_7_9),

    .valid_i_gather_pe              (gather_valid_i_7_9),
    .data_i_gather_pe               (gather_data_i_7_9),
    .ready_o_gather_pe              (gather_ready_o_7_9),
    .valid_o_gather_pe              (gather_valid_o_7_9),
    .data_o_gather_pe               (gather_data_o_7_9),
    .ready_i_gather_pe              (gather_ready_i_7_9),

    .credit_upd                     (credit_upd[7][9])
);


network_interface #(
    .cast_out                       (cast_out_7_10),
    .gather_out                     (gather_out_7_10),
    .cast_sid                       (cast_sid_7_10),
    .gather_sid                     (gather_sid_7_10)
)ni_7_10(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[7][10]),
    .data_i_cast_nw                 (data_o_cast_nw[7][10]),
    .ready_o_cast_nw                (ready_i_cast_nw[7][10]),
    .valid_o_cast_nw                (valid_i_cast_nw[7][10]),
    .data_o_cast_nw                 (data_i_cast_nw[7][10]),
    .ready_i_cast_nw                (ready_o_cast_nw[7][10]),

    .valid_i_gather_nw              (valid_o_gather_nw[7][10]),
    .data_i_gather_nw               (data_o_gather_nw[7][10]),
    .ready_o_gather_nw              (ready_i_gather_nw[7][10]),
    .valid_o_gather_nw              (valid_i_gather_nw[7][10]),
    .data_o_gather_nw               (data_i_gather_nw[7][10]),
    .ready_i_gather_nw              (ready_o_gather_nw[7][10]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[7][10]),
    .data_i_merge_nw                (data_o_merge_nw[7][10]),
    .ready_o_merge_nw               (ready_i_merge_nw[7][10]),
    .valid_o_merge_nw               (valid_i_merge_nw[7][10]),
    .data_o_merge_nw                (data_i_merge_nw[7][10]),
    .ready_i_merge_nw               (ready_o_merge_nw[7][10]),

    .valid_i_cast_pe                (cast_valid_i_7_10),
    .data_i_cast_pe                 (cast_data_i_7_10),
    .ready_o_cast_pe                (cast_ready_o_7_10),
    .valid_o_cast_pe                (cast_valid_o_7_10),
    .data_o_cast_pe                 (cast_data_o_7_10),
    .ready_i_cast_pe                (cast_ready_i_7_10),

    .valid_i_merge_pe               (merge_valid_i_7_10),
    .data_i_merge_pe                (merge_data_i_7_10),
    .ready_o_merge_pe               (merge_ready_o_7_10),
    .valid_o_merge_pe               (merge_valid_o_7_10),
    .data_o_merge_pe                (merge_data_o_7_10),
    .ready_i_merge_pe               (merge_ready_i_7_10),

    .valid_i_gather_pe              (gather_valid_i_7_10),
    .data_i_gather_pe               (gather_data_i_7_10),
    .ready_o_gather_pe              (gather_ready_o_7_10),
    .valid_o_gather_pe              (gather_valid_o_7_10),
    .data_o_gather_pe               (gather_data_o_7_10),
    .ready_i_gather_pe              (gather_ready_i_7_10),

    .credit_upd                     (credit_upd[7][10])
);


network_interface #(
    .cast_out                       (cast_out_7_11),
    .gather_out                     (gather_out_7_11),
    .cast_sid                       (cast_sid_7_11),
    .gather_sid                     (gather_sid_7_11)
)ni_7_11(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[7][11]),
    .data_i_cast_nw                 (data_o_cast_nw[7][11]),
    .ready_o_cast_nw                (ready_i_cast_nw[7][11]),
    .valid_o_cast_nw                (valid_i_cast_nw[7][11]),
    .data_o_cast_nw                 (data_i_cast_nw[7][11]),
    .ready_i_cast_nw                (ready_o_cast_nw[7][11]),

    .valid_i_gather_nw              (valid_o_gather_nw[7][11]),
    .data_i_gather_nw               (data_o_gather_nw[7][11]),
    .ready_o_gather_nw              (ready_i_gather_nw[7][11]),
    .valid_o_gather_nw              (valid_i_gather_nw[7][11]),
    .data_o_gather_nw               (data_i_gather_nw[7][11]),
    .ready_i_gather_nw              (ready_o_gather_nw[7][11]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[7][11]),
    .data_i_merge_nw                (data_o_merge_nw[7][11]),
    .ready_o_merge_nw               (ready_i_merge_nw[7][11]),
    .valid_o_merge_nw               (valid_i_merge_nw[7][11]),
    .data_o_merge_nw                (data_i_merge_nw[7][11]),
    .ready_i_merge_nw               (ready_o_merge_nw[7][11]),

    .valid_i_cast_pe                (cast_valid_i_7_11),
    .data_i_cast_pe                 (cast_data_i_7_11),
    .ready_o_cast_pe                (cast_ready_o_7_11),
    .valid_o_cast_pe                (cast_valid_o_7_11),
    .data_o_cast_pe                 (cast_data_o_7_11),
    .ready_i_cast_pe                (cast_ready_i_7_11),

    .valid_i_merge_pe               (merge_valid_i_7_11),
    .data_i_merge_pe                (merge_data_i_7_11),
    .ready_o_merge_pe               (merge_ready_o_7_11),
    .valid_o_merge_pe               (merge_valid_o_7_11),
    .data_o_merge_pe                (merge_data_o_7_11),
    .ready_i_merge_pe               (merge_ready_i_7_11),

    .valid_i_gather_pe              (gather_valid_i_7_11),
    .data_i_gather_pe               (gather_data_i_7_11),
    .ready_o_gather_pe              (gather_ready_o_7_11),
    .valid_o_gather_pe              (gather_valid_o_7_11),
    .data_o_gather_pe               (gather_data_o_7_11),
    .ready_i_gather_pe              (gather_ready_i_7_11),

    .credit_upd                     (credit_upd[7][11])
);


network_interface #(
    .cast_out                       (cast_out_7_12),
    .gather_out                     (gather_out_7_12),
    .cast_sid                       (cast_sid_7_12),
    .gather_sid                     (gather_sid_7_12)
)ni_7_12(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[7][12]),
    .data_i_cast_nw                 (data_o_cast_nw[7][12]),
    .ready_o_cast_nw                (ready_i_cast_nw[7][12]),
    .valid_o_cast_nw                (valid_i_cast_nw[7][12]),
    .data_o_cast_nw                 (data_i_cast_nw[7][12]),
    .ready_i_cast_nw                (ready_o_cast_nw[7][12]),

    .valid_i_gather_nw              (valid_o_gather_nw[7][12]),
    .data_i_gather_nw               (data_o_gather_nw[7][12]),
    .ready_o_gather_nw              (ready_i_gather_nw[7][12]),
    .valid_o_gather_nw              (valid_i_gather_nw[7][12]),
    .data_o_gather_nw               (data_i_gather_nw[7][12]),
    .ready_i_gather_nw              (ready_o_gather_nw[7][12]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[7][12]),
    .data_i_merge_nw                (data_o_merge_nw[7][12]),
    .ready_o_merge_nw               (ready_i_merge_nw[7][12]),
    .valid_o_merge_nw               (valid_i_merge_nw[7][12]),
    .data_o_merge_nw                (data_i_merge_nw[7][12]),
    .ready_i_merge_nw               (ready_o_merge_nw[7][12]),

    .valid_i_cast_pe                (cast_valid_i_7_12),
    .data_i_cast_pe                 (cast_data_i_7_12),
    .ready_o_cast_pe                (cast_ready_o_7_12),
    .valid_o_cast_pe                (cast_valid_o_7_12),
    .data_o_cast_pe                 (cast_data_o_7_12),
    .ready_i_cast_pe                (cast_ready_i_7_12),

    .valid_i_merge_pe               (merge_valid_i_7_12),
    .data_i_merge_pe                (merge_data_i_7_12),
    .ready_o_merge_pe               (merge_ready_o_7_12),
    .valid_o_merge_pe               (merge_valid_o_7_12),
    .data_o_merge_pe                (merge_data_o_7_12),
    .ready_i_merge_pe               (merge_ready_i_7_12),

    .valid_i_gather_pe              (gather_valid_i_7_12),
    .data_i_gather_pe               (gather_data_i_7_12),
    .ready_o_gather_pe              (gather_ready_o_7_12),
    .valid_o_gather_pe              (gather_valid_o_7_12),
    .data_o_gather_pe               (gather_data_o_7_12),
    .ready_i_gather_pe              (gather_ready_i_7_12),

    .credit_upd                     (credit_upd[7][12])
);


network_interface #(
    .cast_out                       (cast_out_7_13),
    .gather_out                     (gather_out_7_13),
    .cast_sid                       (cast_sid_7_13),
    .gather_sid                     (gather_sid_7_13)
)ni_7_13(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[7][13]),
    .data_i_cast_nw                 (data_o_cast_nw[7][13]),
    .ready_o_cast_nw                (ready_i_cast_nw[7][13]),
    .valid_o_cast_nw                (valid_i_cast_nw[7][13]),
    .data_o_cast_nw                 (data_i_cast_nw[7][13]),
    .ready_i_cast_nw                (ready_o_cast_nw[7][13]),

    .valid_i_gather_nw              (valid_o_gather_nw[7][13]),
    .data_i_gather_nw               (data_o_gather_nw[7][13]),
    .ready_o_gather_nw              (ready_i_gather_nw[7][13]),
    .valid_o_gather_nw              (valid_i_gather_nw[7][13]),
    .data_o_gather_nw               (data_i_gather_nw[7][13]),
    .ready_i_gather_nw              (ready_o_gather_nw[7][13]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[7][13]),
    .data_i_merge_nw                (data_o_merge_nw[7][13]),
    .ready_o_merge_nw               (ready_i_merge_nw[7][13]),
    .valid_o_merge_nw               (valid_i_merge_nw[7][13]),
    .data_o_merge_nw                (data_i_merge_nw[7][13]),
    .ready_i_merge_nw               (ready_o_merge_nw[7][13]),

    .valid_i_cast_pe                (cast_valid_i_7_13),
    .data_i_cast_pe                 (cast_data_i_7_13),
    .ready_o_cast_pe                (cast_ready_o_7_13),
    .valid_o_cast_pe                (cast_valid_o_7_13),
    .data_o_cast_pe                 (cast_data_o_7_13),
    .ready_i_cast_pe                (cast_ready_i_7_13),

    .valid_i_merge_pe               (merge_valid_i_7_13),
    .data_i_merge_pe                (merge_data_i_7_13),
    .ready_o_merge_pe               (merge_ready_o_7_13),
    .valid_o_merge_pe               (merge_valid_o_7_13),
    .data_o_merge_pe                (merge_data_o_7_13),
    .ready_i_merge_pe               (merge_ready_i_7_13),

    .valid_i_gather_pe              (gather_valid_i_7_13),
    .data_i_gather_pe               (gather_data_i_7_13),
    .ready_o_gather_pe              (gather_ready_o_7_13),
    .valid_o_gather_pe              (gather_valid_o_7_13),
    .data_o_gather_pe               (gather_data_o_7_13),
    .ready_i_gather_pe              (gather_ready_i_7_13),

    .credit_upd                     (credit_upd[7][13])
);


network_interface #(
    .cast_out                       (cast_out_7_14),
    .gather_out                     (gather_out_7_14),
    .cast_sid                       (cast_sid_7_14),
    .gather_sid                     (gather_sid_7_14)
)ni_7_14(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[7][14]),
    .data_i_cast_nw                 (data_o_cast_nw[7][14]),
    .ready_o_cast_nw                (ready_i_cast_nw[7][14]),
    .valid_o_cast_nw                (valid_i_cast_nw[7][14]),
    .data_o_cast_nw                 (data_i_cast_nw[7][14]),
    .ready_i_cast_nw                (ready_o_cast_nw[7][14]),

    .valid_i_gather_nw              (valid_o_gather_nw[7][14]),
    .data_i_gather_nw               (data_o_gather_nw[7][14]),
    .ready_o_gather_nw              (ready_i_gather_nw[7][14]),
    .valid_o_gather_nw              (valid_i_gather_nw[7][14]),
    .data_o_gather_nw               (data_i_gather_nw[7][14]),
    .ready_i_gather_nw              (ready_o_gather_nw[7][14]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[7][14]),
    .data_i_merge_nw                (data_o_merge_nw[7][14]),
    .ready_o_merge_nw               (ready_i_merge_nw[7][14]),
    .valid_o_merge_nw               (valid_i_merge_nw[7][14]),
    .data_o_merge_nw                (data_i_merge_nw[7][14]),
    .ready_i_merge_nw               (ready_o_merge_nw[7][14]),

    .valid_i_cast_pe                (cast_valid_i_7_14),
    .data_i_cast_pe                 (cast_data_i_7_14),
    .ready_o_cast_pe                (cast_ready_o_7_14),
    .valid_o_cast_pe                (cast_valid_o_7_14),
    .data_o_cast_pe                 (cast_data_o_7_14),
    .ready_i_cast_pe                (cast_ready_i_7_14),

    .valid_i_merge_pe               (merge_valid_i_7_14),
    .data_i_merge_pe                (merge_data_i_7_14),
    .ready_o_merge_pe               (merge_ready_o_7_14),
    .valid_o_merge_pe               (merge_valid_o_7_14),
    .data_o_merge_pe                (merge_data_o_7_14),
    .ready_i_merge_pe               (merge_ready_i_7_14),

    .valid_i_gather_pe              (gather_valid_i_7_14),
    .data_i_gather_pe               (gather_data_i_7_14),
    .ready_o_gather_pe              (gather_ready_o_7_14),
    .valid_o_gather_pe              (gather_valid_o_7_14),
    .data_o_gather_pe               (gather_data_o_7_14),
    .ready_i_gather_pe              (gather_ready_i_7_14),

    .credit_upd                     (credit_upd[7][14])
);


network_interface #(
    .cast_out                       (cast_out_7_15),
    .gather_out                     (gather_out_7_15),
    .cast_sid                       (cast_sid_7_15),
    .gather_sid                     (gather_sid_7_15)
)ni_7_15(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[7][15]),
    .data_i_cast_nw                 (data_o_cast_nw[7][15]),
    .ready_o_cast_nw                (ready_i_cast_nw[7][15]),
    .valid_o_cast_nw                (valid_i_cast_nw[7][15]),
    .data_o_cast_nw                 (data_i_cast_nw[7][15]),
    .ready_i_cast_nw                (ready_o_cast_nw[7][15]),

    .valid_i_gather_nw              (valid_o_gather_nw[7][15]),
    .data_i_gather_nw               (data_o_gather_nw[7][15]),
    .ready_o_gather_nw              (ready_i_gather_nw[7][15]),
    .valid_o_gather_nw              (valid_i_gather_nw[7][15]),
    .data_o_gather_nw               (data_i_gather_nw[7][15]),
    .ready_i_gather_nw              (ready_o_gather_nw[7][15]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[7][15]),
    .data_i_merge_nw                (data_o_merge_nw[7][15]),
    .ready_o_merge_nw               (ready_i_merge_nw[7][15]),
    .valid_o_merge_nw               (valid_i_merge_nw[7][15]),
    .data_o_merge_nw                (data_i_merge_nw[7][15]),
    .ready_i_merge_nw               (ready_o_merge_nw[7][15]),

    .valid_i_cast_pe                (cast_valid_i_7_15),
    .data_i_cast_pe                 (cast_data_i_7_15),
    .ready_o_cast_pe                (cast_ready_o_7_15),
    .valid_o_cast_pe                (cast_valid_o_7_15),
    .data_o_cast_pe                 (cast_data_o_7_15),
    .ready_i_cast_pe                (cast_ready_i_7_15),

    .valid_i_merge_pe               (merge_valid_i_7_15),
    .data_i_merge_pe                (merge_data_i_7_15),
    .ready_o_merge_pe               (merge_ready_o_7_15),
    .valid_o_merge_pe               (merge_valid_o_7_15),
    .data_o_merge_pe                (merge_data_o_7_15),
    .ready_i_merge_pe               (merge_ready_i_7_15),

    .valid_i_gather_pe              (gather_valid_i_7_15),
    .data_i_gather_pe               (gather_data_i_7_15),
    .ready_o_gather_pe              (gather_ready_o_7_15),
    .valid_o_gather_pe              (gather_valid_o_7_15),
    .data_o_gather_pe               (gather_data_o_7_15),
    .ready_i_gather_pe              (gather_ready_i_7_15),

    .credit_upd                     (credit_upd[7][15])
);


network_interface #(
    .cast_out                       (cast_out_7_16),
    .gather_out                     (gather_out_7_16),
    .cast_sid                       (cast_sid_7_16),
    .gather_sid                     (gather_sid_7_16)
)ni_7_16(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[7][16]),
    .data_i_cast_nw                 (data_o_cast_nw[7][16]),
    .ready_o_cast_nw                (ready_i_cast_nw[7][16]),
    .valid_o_cast_nw                (valid_i_cast_nw[7][16]),
    .data_o_cast_nw                 (data_i_cast_nw[7][16]),
    .ready_i_cast_nw                (ready_o_cast_nw[7][16]),

    .valid_i_gather_nw              (valid_o_gather_nw[7][16]),
    .data_i_gather_nw               (data_o_gather_nw[7][16]),
    .ready_o_gather_nw              (ready_i_gather_nw[7][16]),
    .valid_o_gather_nw              (valid_i_gather_nw[7][16]),
    .data_o_gather_nw               (data_i_gather_nw[7][16]),
    .ready_i_gather_nw              (ready_o_gather_nw[7][16]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[7][16]),
    .data_i_merge_nw                (data_o_merge_nw[7][16]),
    .ready_o_merge_nw               (ready_i_merge_nw[7][16]),
    .valid_o_merge_nw               (valid_i_merge_nw[7][16]),
    .data_o_merge_nw                (data_i_merge_nw[7][16]),
    .ready_i_merge_nw               (ready_o_merge_nw[7][16]),

    .valid_i_cast_pe                (cast_valid_i_7_16),
    .data_i_cast_pe                 (cast_data_i_7_16),
    .ready_o_cast_pe                (cast_ready_o_7_16),
    .valid_o_cast_pe                (cast_valid_o_7_16),
    .data_o_cast_pe                 (cast_data_o_7_16),
    .ready_i_cast_pe                (cast_ready_i_7_16),

    .valid_i_merge_pe               (merge_valid_i_7_16),
    .data_i_merge_pe                (merge_data_i_7_16),
    .ready_o_merge_pe               (merge_ready_o_7_16),
    .valid_o_merge_pe               (merge_valid_o_7_16),
    .data_o_merge_pe                (merge_data_o_7_16),
    .ready_i_merge_pe               (merge_ready_i_7_16),

    .valid_i_gather_pe              (gather_valid_i_7_16),
    .data_i_gather_pe               (gather_data_i_7_16),
    .ready_o_gather_pe              (gather_ready_o_7_16),
    .valid_o_gather_pe              (gather_valid_o_7_16),
    .data_o_gather_pe               (gather_data_o_7_16),
    .ready_i_gather_pe              (gather_ready_i_7_16),

    .credit_upd                     (credit_upd[7][16])
);


network_interface #(
    .cast_out                       (cast_out_7_17),
    .gather_out                     (gather_out_7_17),
    .cast_sid                       (cast_sid_7_17),
    .gather_sid                     (gather_sid_7_17)
)ni_7_17(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[7][17]),
    .data_i_cast_nw                 (data_o_cast_nw[7][17]),
    .ready_o_cast_nw                (ready_i_cast_nw[7][17]),
    .valid_o_cast_nw                (valid_i_cast_nw[7][17]),
    .data_o_cast_nw                 (data_i_cast_nw[7][17]),
    .ready_i_cast_nw                (ready_o_cast_nw[7][17]),

    .valid_i_gather_nw              (valid_o_gather_nw[7][17]),
    .data_i_gather_nw               (data_o_gather_nw[7][17]),
    .ready_o_gather_nw              (ready_i_gather_nw[7][17]),
    .valid_o_gather_nw              (valid_i_gather_nw[7][17]),
    .data_o_gather_nw               (data_i_gather_nw[7][17]),
    .ready_i_gather_nw              (ready_o_gather_nw[7][17]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[7][17]),
    .data_i_merge_nw                (data_o_merge_nw[7][17]),
    .ready_o_merge_nw               (ready_i_merge_nw[7][17]),
    .valid_o_merge_nw               (valid_i_merge_nw[7][17]),
    .data_o_merge_nw                (data_i_merge_nw[7][17]),
    .ready_i_merge_nw               (ready_o_merge_nw[7][17]),

    .valid_i_cast_pe                (cast_valid_i_7_17),
    .data_i_cast_pe                 (cast_data_i_7_17),
    .ready_o_cast_pe                (cast_ready_o_7_17),
    .valid_o_cast_pe                (cast_valid_o_7_17),
    .data_o_cast_pe                 (cast_data_o_7_17),
    .ready_i_cast_pe                (cast_ready_i_7_17),

    .valid_i_merge_pe               (merge_valid_i_7_17),
    .data_i_merge_pe                (merge_data_i_7_17),
    .ready_o_merge_pe               (merge_ready_o_7_17),
    .valid_o_merge_pe               (merge_valid_o_7_17),
    .data_o_merge_pe                (merge_data_o_7_17),
    .ready_i_merge_pe               (merge_ready_i_7_17),

    .valid_i_gather_pe              (gather_valid_i_7_17),
    .data_i_gather_pe               (gather_data_i_7_17),
    .ready_o_gather_pe              (gather_ready_o_7_17),
    .valid_o_gather_pe              (gather_valid_o_7_17),
    .data_o_gather_pe               (gather_data_o_7_17),
    .ready_i_gather_pe              (gather_ready_i_7_17),

    .credit_upd                     (credit_upd[7][17])
);


network_interface #(
    .cast_out                       (cast_out_7_18),
    .gather_out                     (gather_out_7_18),
    .cast_sid                       (cast_sid_7_18),
    .gather_sid                     (gather_sid_7_18)
)ni_7_18(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[7][18]),
    .data_i_cast_nw                 (data_o_cast_nw[7][18]),
    .ready_o_cast_nw                (ready_i_cast_nw[7][18]),
    .valid_o_cast_nw                (valid_i_cast_nw[7][18]),
    .data_o_cast_nw                 (data_i_cast_nw[7][18]),
    .ready_i_cast_nw                (ready_o_cast_nw[7][18]),

    .valid_i_gather_nw              (valid_o_gather_nw[7][18]),
    .data_i_gather_nw               (data_o_gather_nw[7][18]),
    .ready_o_gather_nw              (ready_i_gather_nw[7][18]),
    .valid_o_gather_nw              (valid_i_gather_nw[7][18]),
    .data_o_gather_nw               (data_i_gather_nw[7][18]),
    .ready_i_gather_nw              (ready_o_gather_nw[7][18]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[7][18]),
    .data_i_merge_nw                (data_o_merge_nw[7][18]),
    .ready_o_merge_nw               (ready_i_merge_nw[7][18]),
    .valid_o_merge_nw               (valid_i_merge_nw[7][18]),
    .data_o_merge_nw                (data_i_merge_nw[7][18]),
    .ready_i_merge_nw               (ready_o_merge_nw[7][18]),

    .valid_i_cast_pe                (cast_valid_i_7_18),
    .data_i_cast_pe                 (cast_data_i_7_18),
    .ready_o_cast_pe                (cast_ready_o_7_18),
    .valid_o_cast_pe                (cast_valid_o_7_18),
    .data_o_cast_pe                 (cast_data_o_7_18),
    .ready_i_cast_pe                (cast_ready_i_7_18),

    .valid_i_merge_pe               (merge_valid_i_7_18),
    .data_i_merge_pe                (merge_data_i_7_18),
    .ready_o_merge_pe               (merge_ready_o_7_18),
    .valid_o_merge_pe               (merge_valid_o_7_18),
    .data_o_merge_pe                (merge_data_o_7_18),
    .ready_i_merge_pe               (merge_ready_i_7_18),

    .valid_i_gather_pe              (gather_valid_i_7_18),
    .data_i_gather_pe               (gather_data_i_7_18),
    .ready_o_gather_pe              (gather_ready_o_7_18),
    .valid_o_gather_pe              (gather_valid_o_7_18),
    .data_o_gather_pe               (gather_data_o_7_18),
    .ready_i_gather_pe              (gather_ready_i_7_18),

    .credit_upd                     (credit_upd[7][18])
);


network_interface #(
    .cast_out                       (cast_out_7_19),
    .gather_out                     (gather_out_7_19),
    .cast_sid                       (cast_sid_7_19),
    .gather_sid                     (gather_sid_7_19)
)ni_7_19(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[7][19]),
    .data_i_cast_nw                 (data_o_cast_nw[7][19]),
    .ready_o_cast_nw                (ready_i_cast_nw[7][19]),
    .valid_o_cast_nw                (valid_i_cast_nw[7][19]),
    .data_o_cast_nw                 (data_i_cast_nw[7][19]),
    .ready_i_cast_nw                (ready_o_cast_nw[7][19]),

    .valid_i_gather_nw              (valid_o_gather_nw[7][19]),
    .data_i_gather_nw               (data_o_gather_nw[7][19]),
    .ready_o_gather_nw              (ready_i_gather_nw[7][19]),
    .valid_o_gather_nw              (valid_i_gather_nw[7][19]),
    .data_o_gather_nw               (data_i_gather_nw[7][19]),
    .ready_i_gather_nw              (ready_o_gather_nw[7][19]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[7][19]),
    .data_i_merge_nw                (data_o_merge_nw[7][19]),
    .ready_o_merge_nw               (ready_i_merge_nw[7][19]),
    .valid_o_merge_nw               (valid_i_merge_nw[7][19]),
    .data_o_merge_nw                (data_i_merge_nw[7][19]),
    .ready_i_merge_nw               (ready_o_merge_nw[7][19]),

    .valid_i_cast_pe                (cast_valid_i_7_19),
    .data_i_cast_pe                 (cast_data_i_7_19),
    .ready_o_cast_pe                (cast_ready_o_7_19),
    .valid_o_cast_pe                (cast_valid_o_7_19),
    .data_o_cast_pe                 (cast_data_o_7_19),
    .ready_i_cast_pe                (cast_ready_i_7_19),

    .valid_i_merge_pe               (merge_valid_i_7_19),
    .data_i_merge_pe                (merge_data_i_7_19),
    .ready_o_merge_pe               (merge_ready_o_7_19),
    .valid_o_merge_pe               (merge_valid_o_7_19),
    .data_o_merge_pe                (merge_data_o_7_19),
    .ready_i_merge_pe               (merge_ready_i_7_19),

    .valid_i_gather_pe              (gather_valid_i_7_19),
    .data_i_gather_pe               (gather_data_i_7_19),
    .ready_o_gather_pe              (gather_ready_o_7_19),
    .valid_o_gather_pe              (gather_valid_o_7_19),
    .data_o_gather_pe               (gather_data_o_7_19),
    .ready_i_gather_pe              (gather_ready_i_7_19),

    .credit_upd                     (credit_upd[7][19])
);


network_interface #(
    .cast_out                       (cast_out_7_20),
    .gather_out                     (gather_out_7_20),
    .cast_sid                       (cast_sid_7_20),
    .gather_sid                     (gather_sid_7_20)
)ni_7_20(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[7][20]),
    .data_i_cast_nw                 (data_o_cast_nw[7][20]),
    .ready_o_cast_nw                (ready_i_cast_nw[7][20]),
    .valid_o_cast_nw                (valid_i_cast_nw[7][20]),
    .data_o_cast_nw                 (data_i_cast_nw[7][20]),
    .ready_i_cast_nw                (ready_o_cast_nw[7][20]),

    .valid_i_gather_nw              (valid_o_gather_nw[7][20]),
    .data_i_gather_nw               (data_o_gather_nw[7][20]),
    .ready_o_gather_nw              (ready_i_gather_nw[7][20]),
    .valid_o_gather_nw              (valid_i_gather_nw[7][20]),
    .data_o_gather_nw               (data_i_gather_nw[7][20]),
    .ready_i_gather_nw              (ready_o_gather_nw[7][20]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[7][20]),
    .data_i_merge_nw                (data_o_merge_nw[7][20]),
    .ready_o_merge_nw               (ready_i_merge_nw[7][20]),
    .valid_o_merge_nw               (valid_i_merge_nw[7][20]),
    .data_o_merge_nw                (data_i_merge_nw[7][20]),
    .ready_i_merge_nw               (ready_o_merge_nw[7][20]),

    .valid_i_cast_pe                (cast_valid_i_7_20),
    .data_i_cast_pe                 (cast_data_i_7_20),
    .ready_o_cast_pe                (cast_ready_o_7_20),
    .valid_o_cast_pe                (cast_valid_o_7_20),
    .data_o_cast_pe                 (cast_data_o_7_20),
    .ready_i_cast_pe                (cast_ready_i_7_20),

    .valid_i_merge_pe               (merge_valid_i_7_20),
    .data_i_merge_pe                (merge_data_i_7_20),
    .ready_o_merge_pe               (merge_ready_o_7_20),
    .valid_o_merge_pe               (merge_valid_o_7_20),
    .data_o_merge_pe                (merge_data_o_7_20),
    .ready_i_merge_pe               (merge_ready_i_7_20),

    .valid_i_gather_pe              (gather_valid_i_7_20),
    .data_i_gather_pe               (gather_data_i_7_20),
    .ready_o_gather_pe              (gather_ready_o_7_20),
    .valid_o_gather_pe              (gather_valid_o_7_20),
    .data_o_gather_pe               (gather_data_o_7_20),
    .ready_i_gather_pe              (gather_ready_i_7_20),

    .credit_upd                     (credit_upd[7][20])
);


network_interface #(
    .cast_out                       (cast_out_7_21),
    .gather_out                     (gather_out_7_21),
    .cast_sid                       (cast_sid_7_21),
    .gather_sid                     (gather_sid_7_21)
)ni_7_21(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[7][21]),
    .data_i_cast_nw                 (data_o_cast_nw[7][21]),
    .ready_o_cast_nw                (ready_i_cast_nw[7][21]),
    .valid_o_cast_nw                (valid_i_cast_nw[7][21]),
    .data_o_cast_nw                 (data_i_cast_nw[7][21]),
    .ready_i_cast_nw                (ready_o_cast_nw[7][21]),

    .valid_i_gather_nw              (valid_o_gather_nw[7][21]),
    .data_i_gather_nw               (data_o_gather_nw[7][21]),
    .ready_o_gather_nw              (ready_i_gather_nw[7][21]),
    .valid_o_gather_nw              (valid_i_gather_nw[7][21]),
    .data_o_gather_nw               (data_i_gather_nw[7][21]),
    .ready_i_gather_nw              (ready_o_gather_nw[7][21]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[7][21]),
    .data_i_merge_nw                (data_o_merge_nw[7][21]),
    .ready_o_merge_nw               (ready_i_merge_nw[7][21]),
    .valid_o_merge_nw               (valid_i_merge_nw[7][21]),
    .data_o_merge_nw                (data_i_merge_nw[7][21]),
    .ready_i_merge_nw               (ready_o_merge_nw[7][21]),

    .valid_i_cast_pe                (cast_valid_i_7_21),
    .data_i_cast_pe                 (cast_data_i_7_21),
    .ready_o_cast_pe                (cast_ready_o_7_21),
    .valid_o_cast_pe                (cast_valid_o_7_21),
    .data_o_cast_pe                 (cast_data_o_7_21),
    .ready_i_cast_pe                (cast_ready_i_7_21),

    .valid_i_merge_pe               (merge_valid_i_7_21),
    .data_i_merge_pe                (merge_data_i_7_21),
    .ready_o_merge_pe               (merge_ready_o_7_21),
    .valid_o_merge_pe               (merge_valid_o_7_21),
    .data_o_merge_pe                (merge_data_o_7_21),
    .ready_i_merge_pe               (merge_ready_i_7_21),

    .valid_i_gather_pe              (gather_valid_i_7_21),
    .data_i_gather_pe               (gather_data_i_7_21),
    .ready_o_gather_pe              (gather_ready_o_7_21),
    .valid_o_gather_pe              (gather_valid_o_7_21),
    .data_o_gather_pe               (gather_data_o_7_21),
    .ready_i_gather_pe              (gather_ready_i_7_21),

    .credit_upd                     (credit_upd[7][21])
);


network_interface #(
    .cast_out                       (cast_out_7_22),
    .gather_out                     (gather_out_7_22),
    .cast_sid                       (cast_sid_7_22),
    .gather_sid                     (gather_sid_7_22)
)ni_7_22(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[7][22]),
    .data_i_cast_nw                 (data_o_cast_nw[7][22]),
    .ready_o_cast_nw                (ready_i_cast_nw[7][22]),
    .valid_o_cast_nw                (valid_i_cast_nw[7][22]),
    .data_o_cast_nw                 (data_i_cast_nw[7][22]),
    .ready_i_cast_nw                (ready_o_cast_nw[7][22]),

    .valid_i_gather_nw              (valid_o_gather_nw[7][22]),
    .data_i_gather_nw               (data_o_gather_nw[7][22]),
    .ready_o_gather_nw              (ready_i_gather_nw[7][22]),
    .valid_o_gather_nw              (valid_i_gather_nw[7][22]),
    .data_o_gather_nw               (data_i_gather_nw[7][22]),
    .ready_i_gather_nw              (ready_o_gather_nw[7][22]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[7][22]),
    .data_i_merge_nw                (data_o_merge_nw[7][22]),
    .ready_o_merge_nw               (ready_i_merge_nw[7][22]),
    .valid_o_merge_nw               (valid_i_merge_nw[7][22]),
    .data_o_merge_nw                (data_i_merge_nw[7][22]),
    .ready_i_merge_nw               (ready_o_merge_nw[7][22]),

    .valid_i_cast_pe                (cast_valid_i_7_22),
    .data_i_cast_pe                 (cast_data_i_7_22),
    .ready_o_cast_pe                (cast_ready_o_7_22),
    .valid_o_cast_pe                (cast_valid_o_7_22),
    .data_o_cast_pe                 (cast_data_o_7_22),
    .ready_i_cast_pe                (cast_ready_i_7_22),

    .valid_i_merge_pe               (merge_valid_i_7_22),
    .data_i_merge_pe                (merge_data_i_7_22),
    .ready_o_merge_pe               (merge_ready_o_7_22),
    .valid_o_merge_pe               (merge_valid_o_7_22),
    .data_o_merge_pe                (merge_data_o_7_22),
    .ready_i_merge_pe               (merge_ready_i_7_22),

    .valid_i_gather_pe              (gather_valid_i_7_22),
    .data_i_gather_pe               (gather_data_i_7_22),
    .ready_o_gather_pe              (gather_ready_o_7_22),
    .valid_o_gather_pe              (gather_valid_o_7_22),
    .data_o_gather_pe               (gather_data_o_7_22),
    .ready_i_gather_pe              (gather_ready_i_7_22),

    .credit_upd                     (credit_upd[7][22])
);


network_interface #(
    .cast_out                       (cast_out_7_23),
    .gather_out                     (gather_out_7_23),
    .cast_sid                       (cast_sid_7_23),
    .gather_sid                     (gather_sid_7_23)
)ni_7_23(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[7][23]),
    .data_i_cast_nw                 (data_o_cast_nw[7][23]),
    .ready_o_cast_nw                (ready_i_cast_nw[7][23]),
    .valid_o_cast_nw                (valid_i_cast_nw[7][23]),
    .data_o_cast_nw                 (data_i_cast_nw[7][23]),
    .ready_i_cast_nw                (ready_o_cast_nw[7][23]),

    .valid_i_gather_nw              (valid_o_gather_nw[7][23]),
    .data_i_gather_nw               (data_o_gather_nw[7][23]),
    .ready_o_gather_nw              (ready_i_gather_nw[7][23]),
    .valid_o_gather_nw              (valid_i_gather_nw[7][23]),
    .data_o_gather_nw               (data_i_gather_nw[7][23]),
    .ready_i_gather_nw              (ready_o_gather_nw[7][23]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[7][23]),
    .data_i_merge_nw                (data_o_merge_nw[7][23]),
    .ready_o_merge_nw               (ready_i_merge_nw[7][23]),
    .valid_o_merge_nw               (valid_i_merge_nw[7][23]),
    .data_o_merge_nw                (data_i_merge_nw[7][23]),
    .ready_i_merge_nw               (ready_o_merge_nw[7][23]),

    .valid_i_cast_pe                (cast_valid_i_7_23),
    .data_i_cast_pe                 (cast_data_i_7_23),
    .ready_o_cast_pe                (cast_ready_o_7_23),
    .valid_o_cast_pe                (cast_valid_o_7_23),
    .data_o_cast_pe                 (cast_data_o_7_23),
    .ready_i_cast_pe                (cast_ready_i_7_23),

    .valid_i_merge_pe               (merge_valid_i_7_23),
    .data_i_merge_pe                (merge_data_i_7_23),
    .ready_o_merge_pe               (merge_ready_o_7_23),
    .valid_o_merge_pe               (merge_valid_o_7_23),
    .data_o_merge_pe                (merge_data_o_7_23),
    .ready_i_merge_pe               (merge_ready_i_7_23),

    .valid_i_gather_pe              (gather_valid_i_7_23),
    .data_i_gather_pe               (gather_data_i_7_23),
    .ready_o_gather_pe              (gather_ready_o_7_23),
    .valid_o_gather_pe              (gather_valid_o_7_23),
    .data_o_gather_pe               (gather_data_o_7_23),
    .ready_i_gather_pe              (gather_ready_i_7_23),

    .credit_upd                     (credit_upd[7][23])
);


network_interface #(
    .cast_out                       (cast_out_7_24),
    .gather_out                     (gather_out_7_24),
    .cast_sid                       (cast_sid_7_24),
    .gather_sid                     (gather_sid_7_24)
)ni_7_24(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[7][24]),
    .data_i_cast_nw                 (data_o_cast_nw[7][24]),
    .ready_o_cast_nw                (ready_i_cast_nw[7][24]),
    .valid_o_cast_nw                (valid_i_cast_nw[7][24]),
    .data_o_cast_nw                 (data_i_cast_nw[7][24]),
    .ready_i_cast_nw                (ready_o_cast_nw[7][24]),

    .valid_i_gather_nw              (valid_o_gather_nw[7][24]),
    .data_i_gather_nw               (data_o_gather_nw[7][24]),
    .ready_o_gather_nw              (ready_i_gather_nw[7][24]),
    .valid_o_gather_nw              (valid_i_gather_nw[7][24]),
    .data_o_gather_nw               (data_i_gather_nw[7][24]),
    .ready_i_gather_nw              (ready_o_gather_nw[7][24]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[7][24]),
    .data_i_merge_nw                (data_o_merge_nw[7][24]),
    .ready_o_merge_nw               (ready_i_merge_nw[7][24]),
    .valid_o_merge_nw               (valid_i_merge_nw[7][24]),
    .data_o_merge_nw                (data_i_merge_nw[7][24]),
    .ready_i_merge_nw               (ready_o_merge_nw[7][24]),

    .valid_i_cast_pe                (cast_valid_i_7_24),
    .data_i_cast_pe                 (cast_data_i_7_24),
    .ready_o_cast_pe                (cast_ready_o_7_24),
    .valid_o_cast_pe                (cast_valid_o_7_24),
    .data_o_cast_pe                 (cast_data_o_7_24),
    .ready_i_cast_pe                (cast_ready_i_7_24),

    .valid_i_merge_pe               (merge_valid_i_7_24),
    .data_i_merge_pe                (merge_data_i_7_24),
    .ready_o_merge_pe               (merge_ready_o_7_24),
    .valid_o_merge_pe               (merge_valid_o_7_24),
    .data_o_merge_pe                (merge_data_o_7_24),
    .ready_i_merge_pe               (merge_ready_i_7_24),

    .valid_i_gather_pe              (gather_valid_i_7_24),
    .data_i_gather_pe               (gather_data_i_7_24),
    .ready_o_gather_pe              (gather_ready_o_7_24),
    .valid_o_gather_pe              (gather_valid_o_7_24),
    .data_o_gather_pe               (gather_data_o_7_24),
    .ready_i_gather_pe              (gather_ready_i_7_24),

    .credit_upd                     (credit_upd[7][24])
);


network_interface #(
    .cast_out                       (cast_out_8_0),
    .gather_out                     (gather_out_8_0),
    .cast_sid                       (cast_sid_8_0),
    .gather_sid                     (gather_sid_8_0)
)ni_8_0(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[8][0]),
    .data_i_cast_nw                 (data_o_cast_nw[8][0]),
    .ready_o_cast_nw                (ready_i_cast_nw[8][0]),
    .valid_o_cast_nw                (valid_i_cast_nw[8][0]),
    .data_o_cast_nw                 (data_i_cast_nw[8][0]),
    .ready_i_cast_nw                (ready_o_cast_nw[8][0]),

    .valid_i_gather_nw              (valid_o_gather_nw[8][0]),
    .data_i_gather_nw               (data_o_gather_nw[8][0]),
    .ready_o_gather_nw              (ready_i_gather_nw[8][0]),
    .valid_o_gather_nw              (valid_i_gather_nw[8][0]),
    .data_o_gather_nw               (data_i_gather_nw[8][0]),
    .ready_i_gather_nw              (ready_o_gather_nw[8][0]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[8][0]),
    .data_i_merge_nw                (data_o_merge_nw[8][0]),
    .ready_o_merge_nw               (ready_i_merge_nw[8][0]),
    .valid_o_merge_nw               (valid_i_merge_nw[8][0]),
    .data_o_merge_nw                (data_i_merge_nw[8][0]),
    .ready_i_merge_nw               (ready_o_merge_nw[8][0]),

    .valid_i_cast_pe                (cast_valid_i_8_0),
    .data_i_cast_pe                 (cast_data_i_8_0),
    .ready_o_cast_pe                (cast_ready_o_8_0),
    .valid_o_cast_pe                (cast_valid_o_8_0),
    .data_o_cast_pe                 (cast_data_o_8_0),
    .ready_i_cast_pe                (cast_ready_i_8_0),

    .valid_i_merge_pe               (merge_valid_i_8_0),
    .data_i_merge_pe                (merge_data_i_8_0),
    .ready_o_merge_pe               (merge_ready_o_8_0),
    .valid_o_merge_pe               (merge_valid_o_8_0),
    .data_o_merge_pe                (merge_data_o_8_0),
    .ready_i_merge_pe               (merge_ready_i_8_0),

    .valid_i_gather_pe              (gather_valid_i_8_0),
    .data_i_gather_pe               (gather_data_i_8_0),
    .ready_o_gather_pe              (gather_ready_o_8_0),
    .valid_o_gather_pe              (gather_valid_o_8_0),
    .data_o_gather_pe               (gather_data_o_8_0),
    .ready_i_gather_pe              (gather_ready_i_8_0),

    .credit_upd                     (credit_upd[8][0])
);


network_interface #(
    .cast_out                       (cast_out_8_1),
    .gather_out                     (gather_out_8_1),
    .cast_sid                       (cast_sid_8_1),
    .gather_sid                     (gather_sid_8_1)
)ni_8_1(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[8][1]),
    .data_i_cast_nw                 (data_o_cast_nw[8][1]),
    .ready_o_cast_nw                (ready_i_cast_nw[8][1]),
    .valid_o_cast_nw                (valid_i_cast_nw[8][1]),
    .data_o_cast_nw                 (data_i_cast_nw[8][1]),
    .ready_i_cast_nw                (ready_o_cast_nw[8][1]),

    .valid_i_gather_nw              (valid_o_gather_nw[8][1]),
    .data_i_gather_nw               (data_o_gather_nw[8][1]),
    .ready_o_gather_nw              (ready_i_gather_nw[8][1]),
    .valid_o_gather_nw              (valid_i_gather_nw[8][1]),
    .data_o_gather_nw               (data_i_gather_nw[8][1]),
    .ready_i_gather_nw              (ready_o_gather_nw[8][1]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[8][1]),
    .data_i_merge_nw                (data_o_merge_nw[8][1]),
    .ready_o_merge_nw               (ready_i_merge_nw[8][1]),
    .valid_o_merge_nw               (valid_i_merge_nw[8][1]),
    .data_o_merge_nw                (data_i_merge_nw[8][1]),
    .ready_i_merge_nw               (ready_o_merge_nw[8][1]),

    .valid_i_cast_pe                (cast_valid_i_8_1),
    .data_i_cast_pe                 (cast_data_i_8_1),
    .ready_o_cast_pe                (cast_ready_o_8_1),
    .valid_o_cast_pe                (cast_valid_o_8_1),
    .data_o_cast_pe                 (cast_data_o_8_1),
    .ready_i_cast_pe                (cast_ready_i_8_1),

    .valid_i_merge_pe               (merge_valid_i_8_1),
    .data_i_merge_pe                (merge_data_i_8_1),
    .ready_o_merge_pe               (merge_ready_o_8_1),
    .valid_o_merge_pe               (merge_valid_o_8_1),
    .data_o_merge_pe                (merge_data_o_8_1),
    .ready_i_merge_pe               (merge_ready_i_8_1),

    .valid_i_gather_pe              (gather_valid_i_8_1),
    .data_i_gather_pe               (gather_data_i_8_1),
    .ready_o_gather_pe              (gather_ready_o_8_1),
    .valid_o_gather_pe              (gather_valid_o_8_1),
    .data_o_gather_pe               (gather_data_o_8_1),
    .ready_i_gather_pe              (gather_ready_i_8_1),

    .credit_upd                     (credit_upd[8][1])
);


network_interface #(
    .cast_out                       (cast_out_8_2),
    .gather_out                     (gather_out_8_2),
    .cast_sid                       (cast_sid_8_2),
    .gather_sid                     (gather_sid_8_2)
)ni_8_2(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[8][2]),
    .data_i_cast_nw                 (data_o_cast_nw[8][2]),
    .ready_o_cast_nw                (ready_i_cast_nw[8][2]),
    .valid_o_cast_nw                (valid_i_cast_nw[8][2]),
    .data_o_cast_nw                 (data_i_cast_nw[8][2]),
    .ready_i_cast_nw                (ready_o_cast_nw[8][2]),

    .valid_i_gather_nw              (valid_o_gather_nw[8][2]),
    .data_i_gather_nw               (data_o_gather_nw[8][2]),
    .ready_o_gather_nw              (ready_i_gather_nw[8][2]),
    .valid_o_gather_nw              (valid_i_gather_nw[8][2]),
    .data_o_gather_nw               (data_i_gather_nw[8][2]),
    .ready_i_gather_nw              (ready_o_gather_nw[8][2]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[8][2]),
    .data_i_merge_nw                (data_o_merge_nw[8][2]),
    .ready_o_merge_nw               (ready_i_merge_nw[8][2]),
    .valid_o_merge_nw               (valid_i_merge_nw[8][2]),
    .data_o_merge_nw                (data_i_merge_nw[8][2]),
    .ready_i_merge_nw               (ready_o_merge_nw[8][2]),

    .valid_i_cast_pe                (cast_valid_i_8_2),
    .data_i_cast_pe                 (cast_data_i_8_2),
    .ready_o_cast_pe                (cast_ready_o_8_2),
    .valid_o_cast_pe                (cast_valid_o_8_2),
    .data_o_cast_pe                 (cast_data_o_8_2),
    .ready_i_cast_pe                (cast_ready_i_8_2),

    .valid_i_merge_pe               (merge_valid_i_8_2),
    .data_i_merge_pe                (merge_data_i_8_2),
    .ready_o_merge_pe               (merge_ready_o_8_2),
    .valid_o_merge_pe               (merge_valid_o_8_2),
    .data_o_merge_pe                (merge_data_o_8_2),
    .ready_i_merge_pe               (merge_ready_i_8_2),

    .valid_i_gather_pe              (gather_valid_i_8_2),
    .data_i_gather_pe               (gather_data_i_8_2),
    .ready_o_gather_pe              (gather_ready_o_8_2),
    .valid_o_gather_pe              (gather_valid_o_8_2),
    .data_o_gather_pe               (gather_data_o_8_2),
    .ready_i_gather_pe              (gather_ready_i_8_2),

    .credit_upd                     (credit_upd[8][2])
);


network_interface #(
    .cast_out                       (cast_out_8_3),
    .gather_out                     (gather_out_8_3),
    .cast_sid                       (cast_sid_8_3),
    .gather_sid                     (gather_sid_8_3)
)ni_8_3(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[8][3]),
    .data_i_cast_nw                 (data_o_cast_nw[8][3]),
    .ready_o_cast_nw                (ready_i_cast_nw[8][3]),
    .valid_o_cast_nw                (valid_i_cast_nw[8][3]),
    .data_o_cast_nw                 (data_i_cast_nw[8][3]),
    .ready_i_cast_nw                (ready_o_cast_nw[8][3]),

    .valid_i_gather_nw              (valid_o_gather_nw[8][3]),
    .data_i_gather_nw               (data_o_gather_nw[8][3]),
    .ready_o_gather_nw              (ready_i_gather_nw[8][3]),
    .valid_o_gather_nw              (valid_i_gather_nw[8][3]),
    .data_o_gather_nw               (data_i_gather_nw[8][3]),
    .ready_i_gather_nw              (ready_o_gather_nw[8][3]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[8][3]),
    .data_i_merge_nw                (data_o_merge_nw[8][3]),
    .ready_o_merge_nw               (ready_i_merge_nw[8][3]),
    .valid_o_merge_nw               (valid_i_merge_nw[8][3]),
    .data_o_merge_nw                (data_i_merge_nw[8][3]),
    .ready_i_merge_nw               (ready_o_merge_nw[8][3]),

    .valid_i_cast_pe                (cast_valid_i_8_3),
    .data_i_cast_pe                 (cast_data_i_8_3),
    .ready_o_cast_pe                (cast_ready_o_8_3),
    .valid_o_cast_pe                (cast_valid_o_8_3),
    .data_o_cast_pe                 (cast_data_o_8_3),
    .ready_i_cast_pe                (cast_ready_i_8_3),

    .valid_i_merge_pe               (merge_valid_i_8_3),
    .data_i_merge_pe                (merge_data_i_8_3),
    .ready_o_merge_pe               (merge_ready_o_8_3),
    .valid_o_merge_pe               (merge_valid_o_8_3),
    .data_o_merge_pe                (merge_data_o_8_3),
    .ready_i_merge_pe               (merge_ready_i_8_3),

    .valid_i_gather_pe              (gather_valid_i_8_3),
    .data_i_gather_pe               (gather_data_i_8_3),
    .ready_o_gather_pe              (gather_ready_o_8_3),
    .valid_o_gather_pe              (gather_valid_o_8_3),
    .data_o_gather_pe               (gather_data_o_8_3),
    .ready_i_gather_pe              (gather_ready_i_8_3),

    .credit_upd                     (credit_upd[8][3])
);


network_interface #(
    .cast_out                       (cast_out_8_4),
    .gather_out                     (gather_out_8_4),
    .cast_sid                       (cast_sid_8_4),
    .gather_sid                     (gather_sid_8_4)
)ni_8_4(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[8][4]),
    .data_i_cast_nw                 (data_o_cast_nw[8][4]),
    .ready_o_cast_nw                (ready_i_cast_nw[8][4]),
    .valid_o_cast_nw                (valid_i_cast_nw[8][4]),
    .data_o_cast_nw                 (data_i_cast_nw[8][4]),
    .ready_i_cast_nw                (ready_o_cast_nw[8][4]),

    .valid_i_gather_nw              (valid_o_gather_nw[8][4]),
    .data_i_gather_nw               (data_o_gather_nw[8][4]),
    .ready_o_gather_nw              (ready_i_gather_nw[8][4]),
    .valid_o_gather_nw              (valid_i_gather_nw[8][4]),
    .data_o_gather_nw               (data_i_gather_nw[8][4]),
    .ready_i_gather_nw              (ready_o_gather_nw[8][4]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[8][4]),
    .data_i_merge_nw                (data_o_merge_nw[8][4]),
    .ready_o_merge_nw               (ready_i_merge_nw[8][4]),
    .valid_o_merge_nw               (valid_i_merge_nw[8][4]),
    .data_o_merge_nw                (data_i_merge_nw[8][4]),
    .ready_i_merge_nw               (ready_o_merge_nw[8][4]),

    .valid_i_cast_pe                (cast_valid_i_8_4),
    .data_i_cast_pe                 (cast_data_i_8_4),
    .ready_o_cast_pe                (cast_ready_o_8_4),
    .valid_o_cast_pe                (cast_valid_o_8_4),
    .data_o_cast_pe                 (cast_data_o_8_4),
    .ready_i_cast_pe                (cast_ready_i_8_4),

    .valid_i_merge_pe               (merge_valid_i_8_4),
    .data_i_merge_pe                (merge_data_i_8_4),
    .ready_o_merge_pe               (merge_ready_o_8_4),
    .valid_o_merge_pe               (merge_valid_o_8_4),
    .data_o_merge_pe                (merge_data_o_8_4),
    .ready_i_merge_pe               (merge_ready_i_8_4),

    .valid_i_gather_pe              (gather_valid_i_8_4),
    .data_i_gather_pe               (gather_data_i_8_4),
    .ready_o_gather_pe              (gather_ready_o_8_4),
    .valid_o_gather_pe              (gather_valid_o_8_4),
    .data_o_gather_pe               (gather_data_o_8_4),
    .ready_i_gather_pe              (gather_ready_i_8_4),

    .credit_upd                     (credit_upd[8][4])
);


network_interface #(
    .cast_out                       (cast_out_8_5),
    .gather_out                     (gather_out_8_5),
    .cast_sid                       (cast_sid_8_5),
    .gather_sid                     (gather_sid_8_5)
)ni_8_5(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[8][5]),
    .data_i_cast_nw                 (data_o_cast_nw[8][5]),
    .ready_o_cast_nw                (ready_i_cast_nw[8][5]),
    .valid_o_cast_nw                (valid_i_cast_nw[8][5]),
    .data_o_cast_nw                 (data_i_cast_nw[8][5]),
    .ready_i_cast_nw                (ready_o_cast_nw[8][5]),

    .valid_i_gather_nw              (valid_o_gather_nw[8][5]),
    .data_i_gather_nw               (data_o_gather_nw[8][5]),
    .ready_o_gather_nw              (ready_i_gather_nw[8][5]),
    .valid_o_gather_nw              (valid_i_gather_nw[8][5]),
    .data_o_gather_nw               (data_i_gather_nw[8][5]),
    .ready_i_gather_nw              (ready_o_gather_nw[8][5]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[8][5]),
    .data_i_merge_nw                (data_o_merge_nw[8][5]),
    .ready_o_merge_nw               (ready_i_merge_nw[8][5]),
    .valid_o_merge_nw               (valid_i_merge_nw[8][5]),
    .data_o_merge_nw                (data_i_merge_nw[8][5]),
    .ready_i_merge_nw               (ready_o_merge_nw[8][5]),

    .valid_i_cast_pe                (cast_valid_i_8_5),
    .data_i_cast_pe                 (cast_data_i_8_5),
    .ready_o_cast_pe                (cast_ready_o_8_5),
    .valid_o_cast_pe                (cast_valid_o_8_5),
    .data_o_cast_pe                 (cast_data_o_8_5),
    .ready_i_cast_pe                (cast_ready_i_8_5),

    .valid_i_merge_pe               (merge_valid_i_8_5),
    .data_i_merge_pe                (merge_data_i_8_5),
    .ready_o_merge_pe               (merge_ready_o_8_5),
    .valid_o_merge_pe               (merge_valid_o_8_5),
    .data_o_merge_pe                (merge_data_o_8_5),
    .ready_i_merge_pe               (merge_ready_i_8_5),

    .valid_i_gather_pe              (gather_valid_i_8_5),
    .data_i_gather_pe               (gather_data_i_8_5),
    .ready_o_gather_pe              (gather_ready_o_8_5),
    .valid_o_gather_pe              (gather_valid_o_8_5),
    .data_o_gather_pe               (gather_data_o_8_5),
    .ready_i_gather_pe              (gather_ready_i_8_5),

    .credit_upd                     (credit_upd[8][5])
);


network_interface #(
    .cast_out                       (cast_out_8_6),
    .gather_out                     (gather_out_8_6),
    .cast_sid                       (cast_sid_8_6),
    .gather_sid                     (gather_sid_8_6)
)ni_8_6(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[8][6]),
    .data_i_cast_nw                 (data_o_cast_nw[8][6]),
    .ready_o_cast_nw                (ready_i_cast_nw[8][6]),
    .valid_o_cast_nw                (valid_i_cast_nw[8][6]),
    .data_o_cast_nw                 (data_i_cast_nw[8][6]),
    .ready_i_cast_nw                (ready_o_cast_nw[8][6]),

    .valid_i_gather_nw              (valid_o_gather_nw[8][6]),
    .data_i_gather_nw               (data_o_gather_nw[8][6]),
    .ready_o_gather_nw              (ready_i_gather_nw[8][6]),
    .valid_o_gather_nw              (valid_i_gather_nw[8][6]),
    .data_o_gather_nw               (data_i_gather_nw[8][6]),
    .ready_i_gather_nw              (ready_o_gather_nw[8][6]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[8][6]),
    .data_i_merge_nw                (data_o_merge_nw[8][6]),
    .ready_o_merge_nw               (ready_i_merge_nw[8][6]),
    .valid_o_merge_nw               (valid_i_merge_nw[8][6]),
    .data_o_merge_nw                (data_i_merge_nw[8][6]),
    .ready_i_merge_nw               (ready_o_merge_nw[8][6]),

    .valid_i_cast_pe                (cast_valid_i_8_6),
    .data_i_cast_pe                 (cast_data_i_8_6),
    .ready_o_cast_pe                (cast_ready_o_8_6),
    .valid_o_cast_pe                (cast_valid_o_8_6),
    .data_o_cast_pe                 (cast_data_o_8_6),
    .ready_i_cast_pe                (cast_ready_i_8_6),

    .valid_i_merge_pe               (merge_valid_i_8_6),
    .data_i_merge_pe                (merge_data_i_8_6),
    .ready_o_merge_pe               (merge_ready_o_8_6),
    .valid_o_merge_pe               (merge_valid_o_8_6),
    .data_o_merge_pe                (merge_data_o_8_6),
    .ready_i_merge_pe               (merge_ready_i_8_6),

    .valid_i_gather_pe              (gather_valid_i_8_6),
    .data_i_gather_pe               (gather_data_i_8_6),
    .ready_o_gather_pe              (gather_ready_o_8_6),
    .valid_o_gather_pe              (gather_valid_o_8_6),
    .data_o_gather_pe               (gather_data_o_8_6),
    .ready_i_gather_pe              (gather_ready_i_8_6),

    .credit_upd                     (credit_upd[8][6])
);


network_interface #(
    .cast_out                       (cast_out_8_7),
    .gather_out                     (gather_out_8_7),
    .cast_sid                       (cast_sid_8_7),
    .gather_sid                     (gather_sid_8_7)
)ni_8_7(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[8][7]),
    .data_i_cast_nw                 (data_o_cast_nw[8][7]),
    .ready_o_cast_nw                (ready_i_cast_nw[8][7]),
    .valid_o_cast_nw                (valid_i_cast_nw[8][7]),
    .data_o_cast_nw                 (data_i_cast_nw[8][7]),
    .ready_i_cast_nw                (ready_o_cast_nw[8][7]),

    .valid_i_gather_nw              (valid_o_gather_nw[8][7]),
    .data_i_gather_nw               (data_o_gather_nw[8][7]),
    .ready_o_gather_nw              (ready_i_gather_nw[8][7]),
    .valid_o_gather_nw              (valid_i_gather_nw[8][7]),
    .data_o_gather_nw               (data_i_gather_nw[8][7]),
    .ready_i_gather_nw              (ready_o_gather_nw[8][7]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[8][7]),
    .data_i_merge_nw                (data_o_merge_nw[8][7]),
    .ready_o_merge_nw               (ready_i_merge_nw[8][7]),
    .valid_o_merge_nw               (valid_i_merge_nw[8][7]),
    .data_o_merge_nw                (data_i_merge_nw[8][7]),
    .ready_i_merge_nw               (ready_o_merge_nw[8][7]),

    .valid_i_cast_pe                (cast_valid_i_8_7),
    .data_i_cast_pe                 (cast_data_i_8_7),
    .ready_o_cast_pe                (cast_ready_o_8_7),
    .valid_o_cast_pe                (cast_valid_o_8_7),
    .data_o_cast_pe                 (cast_data_o_8_7),
    .ready_i_cast_pe                (cast_ready_i_8_7),

    .valid_i_merge_pe               (merge_valid_i_8_7),
    .data_i_merge_pe                (merge_data_i_8_7),
    .ready_o_merge_pe               (merge_ready_o_8_7),
    .valid_o_merge_pe               (merge_valid_o_8_7),
    .data_o_merge_pe                (merge_data_o_8_7),
    .ready_i_merge_pe               (merge_ready_i_8_7),

    .valid_i_gather_pe              (gather_valid_i_8_7),
    .data_i_gather_pe               (gather_data_i_8_7),
    .ready_o_gather_pe              (gather_ready_o_8_7),
    .valid_o_gather_pe              (gather_valid_o_8_7),
    .data_o_gather_pe               (gather_data_o_8_7),
    .ready_i_gather_pe              (gather_ready_i_8_7),

    .credit_upd                     (credit_upd[8][7])
);


network_interface #(
    .cast_out                       (cast_out_8_8),
    .gather_out                     (gather_out_8_8),
    .cast_sid                       (cast_sid_8_8),
    .gather_sid                     (gather_sid_8_8)
)ni_8_8(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[8][8]),
    .data_i_cast_nw                 (data_o_cast_nw[8][8]),
    .ready_o_cast_nw                (ready_i_cast_nw[8][8]),
    .valid_o_cast_nw                (valid_i_cast_nw[8][8]),
    .data_o_cast_nw                 (data_i_cast_nw[8][8]),
    .ready_i_cast_nw                (ready_o_cast_nw[8][8]),

    .valid_i_gather_nw              (valid_o_gather_nw[8][8]),
    .data_i_gather_nw               (data_o_gather_nw[8][8]),
    .ready_o_gather_nw              (ready_i_gather_nw[8][8]),
    .valid_o_gather_nw              (valid_i_gather_nw[8][8]),
    .data_o_gather_nw               (data_i_gather_nw[8][8]),
    .ready_i_gather_nw              (ready_o_gather_nw[8][8]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[8][8]),
    .data_i_merge_nw                (data_o_merge_nw[8][8]),
    .ready_o_merge_nw               (ready_i_merge_nw[8][8]),
    .valid_o_merge_nw               (valid_i_merge_nw[8][8]),
    .data_o_merge_nw                (data_i_merge_nw[8][8]),
    .ready_i_merge_nw               (ready_o_merge_nw[8][8]),

    .valid_i_cast_pe                (cast_valid_i_8_8),
    .data_i_cast_pe                 (cast_data_i_8_8),
    .ready_o_cast_pe                (cast_ready_o_8_8),
    .valid_o_cast_pe                (cast_valid_o_8_8),
    .data_o_cast_pe                 (cast_data_o_8_8),
    .ready_i_cast_pe                (cast_ready_i_8_8),

    .valid_i_merge_pe               (merge_valid_i_8_8),
    .data_i_merge_pe                (merge_data_i_8_8),
    .ready_o_merge_pe               (merge_ready_o_8_8),
    .valid_o_merge_pe               (merge_valid_o_8_8),
    .data_o_merge_pe                (merge_data_o_8_8),
    .ready_i_merge_pe               (merge_ready_i_8_8),

    .valid_i_gather_pe              (gather_valid_i_8_8),
    .data_i_gather_pe               (gather_data_i_8_8),
    .ready_o_gather_pe              (gather_ready_o_8_8),
    .valid_o_gather_pe              (gather_valid_o_8_8),
    .data_o_gather_pe               (gather_data_o_8_8),
    .ready_i_gather_pe              (gather_ready_i_8_8),

    .credit_upd                     (credit_upd[8][8])
);


network_interface #(
    .cast_out                       (cast_out_8_9),
    .gather_out                     (gather_out_8_9),
    .cast_sid                       (cast_sid_8_9),
    .gather_sid                     (gather_sid_8_9)
)ni_8_9(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[8][9]),
    .data_i_cast_nw                 (data_o_cast_nw[8][9]),
    .ready_o_cast_nw                (ready_i_cast_nw[8][9]),
    .valid_o_cast_nw                (valid_i_cast_nw[8][9]),
    .data_o_cast_nw                 (data_i_cast_nw[8][9]),
    .ready_i_cast_nw                (ready_o_cast_nw[8][9]),

    .valid_i_gather_nw              (valid_o_gather_nw[8][9]),
    .data_i_gather_nw               (data_o_gather_nw[8][9]),
    .ready_o_gather_nw              (ready_i_gather_nw[8][9]),
    .valid_o_gather_nw              (valid_i_gather_nw[8][9]),
    .data_o_gather_nw               (data_i_gather_nw[8][9]),
    .ready_i_gather_nw              (ready_o_gather_nw[8][9]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[8][9]),
    .data_i_merge_nw                (data_o_merge_nw[8][9]),
    .ready_o_merge_nw               (ready_i_merge_nw[8][9]),
    .valid_o_merge_nw               (valid_i_merge_nw[8][9]),
    .data_o_merge_nw                (data_i_merge_nw[8][9]),
    .ready_i_merge_nw               (ready_o_merge_nw[8][9]),

    .valid_i_cast_pe                (cast_valid_i_8_9),
    .data_i_cast_pe                 (cast_data_i_8_9),
    .ready_o_cast_pe                (cast_ready_o_8_9),
    .valid_o_cast_pe                (cast_valid_o_8_9),
    .data_o_cast_pe                 (cast_data_o_8_9),
    .ready_i_cast_pe                (cast_ready_i_8_9),

    .valid_i_merge_pe               (merge_valid_i_8_9),
    .data_i_merge_pe                (merge_data_i_8_9),
    .ready_o_merge_pe               (merge_ready_o_8_9),
    .valid_o_merge_pe               (merge_valid_o_8_9),
    .data_o_merge_pe                (merge_data_o_8_9),
    .ready_i_merge_pe               (merge_ready_i_8_9),

    .valid_i_gather_pe              (gather_valid_i_8_9),
    .data_i_gather_pe               (gather_data_i_8_9),
    .ready_o_gather_pe              (gather_ready_o_8_9),
    .valid_o_gather_pe              (gather_valid_o_8_9),
    .data_o_gather_pe               (gather_data_o_8_9),
    .ready_i_gather_pe              (gather_ready_i_8_9),

    .credit_upd                     (credit_upd[8][9])
);


network_interface #(
    .cast_out                       (cast_out_8_10),
    .gather_out                     (gather_out_8_10),
    .cast_sid                       (cast_sid_8_10),
    .gather_sid                     (gather_sid_8_10)
)ni_8_10(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[8][10]),
    .data_i_cast_nw                 (data_o_cast_nw[8][10]),
    .ready_o_cast_nw                (ready_i_cast_nw[8][10]),
    .valid_o_cast_nw                (valid_i_cast_nw[8][10]),
    .data_o_cast_nw                 (data_i_cast_nw[8][10]),
    .ready_i_cast_nw                (ready_o_cast_nw[8][10]),

    .valid_i_gather_nw              (valid_o_gather_nw[8][10]),
    .data_i_gather_nw               (data_o_gather_nw[8][10]),
    .ready_o_gather_nw              (ready_i_gather_nw[8][10]),
    .valid_o_gather_nw              (valid_i_gather_nw[8][10]),
    .data_o_gather_nw               (data_i_gather_nw[8][10]),
    .ready_i_gather_nw              (ready_o_gather_nw[8][10]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[8][10]),
    .data_i_merge_nw                (data_o_merge_nw[8][10]),
    .ready_o_merge_nw               (ready_i_merge_nw[8][10]),
    .valid_o_merge_nw               (valid_i_merge_nw[8][10]),
    .data_o_merge_nw                (data_i_merge_nw[8][10]),
    .ready_i_merge_nw               (ready_o_merge_nw[8][10]),

    .valid_i_cast_pe                (cast_valid_i_8_10),
    .data_i_cast_pe                 (cast_data_i_8_10),
    .ready_o_cast_pe                (cast_ready_o_8_10),
    .valid_o_cast_pe                (cast_valid_o_8_10),
    .data_o_cast_pe                 (cast_data_o_8_10),
    .ready_i_cast_pe                (cast_ready_i_8_10),

    .valid_i_merge_pe               (merge_valid_i_8_10),
    .data_i_merge_pe                (merge_data_i_8_10),
    .ready_o_merge_pe               (merge_ready_o_8_10),
    .valid_o_merge_pe               (merge_valid_o_8_10),
    .data_o_merge_pe                (merge_data_o_8_10),
    .ready_i_merge_pe               (merge_ready_i_8_10),

    .valid_i_gather_pe              (gather_valid_i_8_10),
    .data_i_gather_pe               (gather_data_i_8_10),
    .ready_o_gather_pe              (gather_ready_o_8_10),
    .valid_o_gather_pe              (gather_valid_o_8_10),
    .data_o_gather_pe               (gather_data_o_8_10),
    .ready_i_gather_pe              (gather_ready_i_8_10),

    .credit_upd                     (credit_upd[8][10])
);


network_interface #(
    .cast_out                       (cast_out_8_11),
    .gather_out                     (gather_out_8_11),
    .cast_sid                       (cast_sid_8_11),
    .gather_sid                     (gather_sid_8_11)
)ni_8_11(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[8][11]),
    .data_i_cast_nw                 (data_o_cast_nw[8][11]),
    .ready_o_cast_nw                (ready_i_cast_nw[8][11]),
    .valid_o_cast_nw                (valid_i_cast_nw[8][11]),
    .data_o_cast_nw                 (data_i_cast_nw[8][11]),
    .ready_i_cast_nw                (ready_o_cast_nw[8][11]),

    .valid_i_gather_nw              (valid_o_gather_nw[8][11]),
    .data_i_gather_nw               (data_o_gather_nw[8][11]),
    .ready_o_gather_nw              (ready_i_gather_nw[8][11]),
    .valid_o_gather_nw              (valid_i_gather_nw[8][11]),
    .data_o_gather_nw               (data_i_gather_nw[8][11]),
    .ready_i_gather_nw              (ready_o_gather_nw[8][11]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[8][11]),
    .data_i_merge_nw                (data_o_merge_nw[8][11]),
    .ready_o_merge_nw               (ready_i_merge_nw[8][11]),
    .valid_o_merge_nw               (valid_i_merge_nw[8][11]),
    .data_o_merge_nw                (data_i_merge_nw[8][11]),
    .ready_i_merge_nw               (ready_o_merge_nw[8][11]),

    .valid_i_cast_pe                (cast_valid_i_8_11),
    .data_i_cast_pe                 (cast_data_i_8_11),
    .ready_o_cast_pe                (cast_ready_o_8_11),
    .valid_o_cast_pe                (cast_valid_o_8_11),
    .data_o_cast_pe                 (cast_data_o_8_11),
    .ready_i_cast_pe                (cast_ready_i_8_11),

    .valid_i_merge_pe               (merge_valid_i_8_11),
    .data_i_merge_pe                (merge_data_i_8_11),
    .ready_o_merge_pe               (merge_ready_o_8_11),
    .valid_o_merge_pe               (merge_valid_o_8_11),
    .data_o_merge_pe                (merge_data_o_8_11),
    .ready_i_merge_pe               (merge_ready_i_8_11),

    .valid_i_gather_pe              (gather_valid_i_8_11),
    .data_i_gather_pe               (gather_data_i_8_11),
    .ready_o_gather_pe              (gather_ready_o_8_11),
    .valid_o_gather_pe              (gather_valid_o_8_11),
    .data_o_gather_pe               (gather_data_o_8_11),
    .ready_i_gather_pe              (gather_ready_i_8_11),

    .credit_upd                     (credit_upd[8][11])
);


network_interface #(
    .cast_out                       (cast_out_8_12),
    .gather_out                     (gather_out_8_12),
    .cast_sid                       (cast_sid_8_12),
    .gather_sid                     (gather_sid_8_12)
)ni_8_12(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[8][12]),
    .data_i_cast_nw                 (data_o_cast_nw[8][12]),
    .ready_o_cast_nw                (ready_i_cast_nw[8][12]),
    .valid_o_cast_nw                (valid_i_cast_nw[8][12]),
    .data_o_cast_nw                 (data_i_cast_nw[8][12]),
    .ready_i_cast_nw                (ready_o_cast_nw[8][12]),

    .valid_i_gather_nw              (valid_o_gather_nw[8][12]),
    .data_i_gather_nw               (data_o_gather_nw[8][12]),
    .ready_o_gather_nw              (ready_i_gather_nw[8][12]),
    .valid_o_gather_nw              (valid_i_gather_nw[8][12]),
    .data_o_gather_nw               (data_i_gather_nw[8][12]),
    .ready_i_gather_nw              (ready_o_gather_nw[8][12]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[8][12]),
    .data_i_merge_nw                (data_o_merge_nw[8][12]),
    .ready_o_merge_nw               (ready_i_merge_nw[8][12]),
    .valid_o_merge_nw               (valid_i_merge_nw[8][12]),
    .data_o_merge_nw                (data_i_merge_nw[8][12]),
    .ready_i_merge_nw               (ready_o_merge_nw[8][12]),

    .valid_i_cast_pe                (cast_valid_i_8_12),
    .data_i_cast_pe                 (cast_data_i_8_12),
    .ready_o_cast_pe                (cast_ready_o_8_12),
    .valid_o_cast_pe                (cast_valid_o_8_12),
    .data_o_cast_pe                 (cast_data_o_8_12),
    .ready_i_cast_pe                (cast_ready_i_8_12),

    .valid_i_merge_pe               (merge_valid_i_8_12),
    .data_i_merge_pe                (merge_data_i_8_12),
    .ready_o_merge_pe               (merge_ready_o_8_12),
    .valid_o_merge_pe               (merge_valid_o_8_12),
    .data_o_merge_pe                (merge_data_o_8_12),
    .ready_i_merge_pe               (merge_ready_i_8_12),

    .valid_i_gather_pe              (gather_valid_i_8_12),
    .data_i_gather_pe               (gather_data_i_8_12),
    .ready_o_gather_pe              (gather_ready_o_8_12),
    .valid_o_gather_pe              (gather_valid_o_8_12),
    .data_o_gather_pe               (gather_data_o_8_12),
    .ready_i_gather_pe              (gather_ready_i_8_12),

    .credit_upd                     (credit_upd[8][12])
);


network_interface #(
    .cast_out                       (cast_out_8_13),
    .gather_out                     (gather_out_8_13),
    .cast_sid                       (cast_sid_8_13),
    .gather_sid                     (gather_sid_8_13)
)ni_8_13(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[8][13]),
    .data_i_cast_nw                 (data_o_cast_nw[8][13]),
    .ready_o_cast_nw                (ready_i_cast_nw[8][13]),
    .valid_o_cast_nw                (valid_i_cast_nw[8][13]),
    .data_o_cast_nw                 (data_i_cast_nw[8][13]),
    .ready_i_cast_nw                (ready_o_cast_nw[8][13]),

    .valid_i_gather_nw              (valid_o_gather_nw[8][13]),
    .data_i_gather_nw               (data_o_gather_nw[8][13]),
    .ready_o_gather_nw              (ready_i_gather_nw[8][13]),
    .valid_o_gather_nw              (valid_i_gather_nw[8][13]),
    .data_o_gather_nw               (data_i_gather_nw[8][13]),
    .ready_i_gather_nw              (ready_o_gather_nw[8][13]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[8][13]),
    .data_i_merge_nw                (data_o_merge_nw[8][13]),
    .ready_o_merge_nw               (ready_i_merge_nw[8][13]),
    .valid_o_merge_nw               (valid_i_merge_nw[8][13]),
    .data_o_merge_nw                (data_i_merge_nw[8][13]),
    .ready_i_merge_nw               (ready_o_merge_nw[8][13]),

    .valid_i_cast_pe                (cast_valid_i_8_13),
    .data_i_cast_pe                 (cast_data_i_8_13),
    .ready_o_cast_pe                (cast_ready_o_8_13),
    .valid_o_cast_pe                (cast_valid_o_8_13),
    .data_o_cast_pe                 (cast_data_o_8_13),
    .ready_i_cast_pe                (cast_ready_i_8_13),

    .valid_i_merge_pe               (merge_valid_i_8_13),
    .data_i_merge_pe                (merge_data_i_8_13),
    .ready_o_merge_pe               (merge_ready_o_8_13),
    .valid_o_merge_pe               (merge_valid_o_8_13),
    .data_o_merge_pe                (merge_data_o_8_13),
    .ready_i_merge_pe               (merge_ready_i_8_13),

    .valid_i_gather_pe              (gather_valid_i_8_13),
    .data_i_gather_pe               (gather_data_i_8_13),
    .ready_o_gather_pe              (gather_ready_o_8_13),
    .valid_o_gather_pe              (gather_valid_o_8_13),
    .data_o_gather_pe               (gather_data_o_8_13),
    .ready_i_gather_pe              (gather_ready_i_8_13),

    .credit_upd                     (credit_upd[8][13])
);


network_interface #(
    .cast_out                       (cast_out_8_14),
    .gather_out                     (gather_out_8_14),
    .cast_sid                       (cast_sid_8_14),
    .gather_sid                     (gather_sid_8_14)
)ni_8_14(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[8][14]),
    .data_i_cast_nw                 (data_o_cast_nw[8][14]),
    .ready_o_cast_nw                (ready_i_cast_nw[8][14]),
    .valid_o_cast_nw                (valid_i_cast_nw[8][14]),
    .data_o_cast_nw                 (data_i_cast_nw[8][14]),
    .ready_i_cast_nw                (ready_o_cast_nw[8][14]),

    .valid_i_gather_nw              (valid_o_gather_nw[8][14]),
    .data_i_gather_nw               (data_o_gather_nw[8][14]),
    .ready_o_gather_nw              (ready_i_gather_nw[8][14]),
    .valid_o_gather_nw              (valid_i_gather_nw[8][14]),
    .data_o_gather_nw               (data_i_gather_nw[8][14]),
    .ready_i_gather_nw              (ready_o_gather_nw[8][14]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[8][14]),
    .data_i_merge_nw                (data_o_merge_nw[8][14]),
    .ready_o_merge_nw               (ready_i_merge_nw[8][14]),
    .valid_o_merge_nw               (valid_i_merge_nw[8][14]),
    .data_o_merge_nw                (data_i_merge_nw[8][14]),
    .ready_i_merge_nw               (ready_o_merge_nw[8][14]),

    .valid_i_cast_pe                (cast_valid_i_8_14),
    .data_i_cast_pe                 (cast_data_i_8_14),
    .ready_o_cast_pe                (cast_ready_o_8_14),
    .valid_o_cast_pe                (cast_valid_o_8_14),
    .data_o_cast_pe                 (cast_data_o_8_14),
    .ready_i_cast_pe                (cast_ready_i_8_14),

    .valid_i_merge_pe               (merge_valid_i_8_14),
    .data_i_merge_pe                (merge_data_i_8_14),
    .ready_o_merge_pe               (merge_ready_o_8_14),
    .valid_o_merge_pe               (merge_valid_o_8_14),
    .data_o_merge_pe                (merge_data_o_8_14),
    .ready_i_merge_pe               (merge_ready_i_8_14),

    .valid_i_gather_pe              (gather_valid_i_8_14),
    .data_i_gather_pe               (gather_data_i_8_14),
    .ready_o_gather_pe              (gather_ready_o_8_14),
    .valid_o_gather_pe              (gather_valid_o_8_14),
    .data_o_gather_pe               (gather_data_o_8_14),
    .ready_i_gather_pe              (gather_ready_i_8_14),

    .credit_upd                     (credit_upd[8][14])
);


network_interface #(
    .cast_out                       (cast_out_8_15),
    .gather_out                     (gather_out_8_15),
    .cast_sid                       (cast_sid_8_15),
    .gather_sid                     (gather_sid_8_15)
)ni_8_15(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[8][15]),
    .data_i_cast_nw                 (data_o_cast_nw[8][15]),
    .ready_o_cast_nw                (ready_i_cast_nw[8][15]),
    .valid_o_cast_nw                (valid_i_cast_nw[8][15]),
    .data_o_cast_nw                 (data_i_cast_nw[8][15]),
    .ready_i_cast_nw                (ready_o_cast_nw[8][15]),

    .valid_i_gather_nw              (valid_o_gather_nw[8][15]),
    .data_i_gather_nw               (data_o_gather_nw[8][15]),
    .ready_o_gather_nw              (ready_i_gather_nw[8][15]),
    .valid_o_gather_nw              (valid_i_gather_nw[8][15]),
    .data_o_gather_nw               (data_i_gather_nw[8][15]),
    .ready_i_gather_nw              (ready_o_gather_nw[8][15]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[8][15]),
    .data_i_merge_nw                (data_o_merge_nw[8][15]),
    .ready_o_merge_nw               (ready_i_merge_nw[8][15]),
    .valid_o_merge_nw               (valid_i_merge_nw[8][15]),
    .data_o_merge_nw                (data_i_merge_nw[8][15]),
    .ready_i_merge_nw               (ready_o_merge_nw[8][15]),

    .valid_i_cast_pe                (cast_valid_i_8_15),
    .data_i_cast_pe                 (cast_data_i_8_15),
    .ready_o_cast_pe                (cast_ready_o_8_15),
    .valid_o_cast_pe                (cast_valid_o_8_15),
    .data_o_cast_pe                 (cast_data_o_8_15),
    .ready_i_cast_pe                (cast_ready_i_8_15),

    .valid_i_merge_pe               (merge_valid_i_8_15),
    .data_i_merge_pe                (merge_data_i_8_15),
    .ready_o_merge_pe               (merge_ready_o_8_15),
    .valid_o_merge_pe               (merge_valid_o_8_15),
    .data_o_merge_pe                (merge_data_o_8_15),
    .ready_i_merge_pe               (merge_ready_i_8_15),

    .valid_i_gather_pe              (gather_valid_i_8_15),
    .data_i_gather_pe               (gather_data_i_8_15),
    .ready_o_gather_pe              (gather_ready_o_8_15),
    .valid_o_gather_pe              (gather_valid_o_8_15),
    .data_o_gather_pe               (gather_data_o_8_15),
    .ready_i_gather_pe              (gather_ready_i_8_15),

    .credit_upd                     (credit_upd[8][15])
);


network_interface #(
    .cast_out                       (cast_out_8_16),
    .gather_out                     (gather_out_8_16),
    .cast_sid                       (cast_sid_8_16),
    .gather_sid                     (gather_sid_8_16)
)ni_8_16(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[8][16]),
    .data_i_cast_nw                 (data_o_cast_nw[8][16]),
    .ready_o_cast_nw                (ready_i_cast_nw[8][16]),
    .valid_o_cast_nw                (valid_i_cast_nw[8][16]),
    .data_o_cast_nw                 (data_i_cast_nw[8][16]),
    .ready_i_cast_nw                (ready_o_cast_nw[8][16]),

    .valid_i_gather_nw              (valid_o_gather_nw[8][16]),
    .data_i_gather_nw               (data_o_gather_nw[8][16]),
    .ready_o_gather_nw              (ready_i_gather_nw[8][16]),
    .valid_o_gather_nw              (valid_i_gather_nw[8][16]),
    .data_o_gather_nw               (data_i_gather_nw[8][16]),
    .ready_i_gather_nw              (ready_o_gather_nw[8][16]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[8][16]),
    .data_i_merge_nw                (data_o_merge_nw[8][16]),
    .ready_o_merge_nw               (ready_i_merge_nw[8][16]),
    .valid_o_merge_nw               (valid_i_merge_nw[8][16]),
    .data_o_merge_nw                (data_i_merge_nw[8][16]),
    .ready_i_merge_nw               (ready_o_merge_nw[8][16]),

    .valid_i_cast_pe                (cast_valid_i_8_16),
    .data_i_cast_pe                 (cast_data_i_8_16),
    .ready_o_cast_pe                (cast_ready_o_8_16),
    .valid_o_cast_pe                (cast_valid_o_8_16),
    .data_o_cast_pe                 (cast_data_o_8_16),
    .ready_i_cast_pe                (cast_ready_i_8_16),

    .valid_i_merge_pe               (merge_valid_i_8_16),
    .data_i_merge_pe                (merge_data_i_8_16),
    .ready_o_merge_pe               (merge_ready_o_8_16),
    .valid_o_merge_pe               (merge_valid_o_8_16),
    .data_o_merge_pe                (merge_data_o_8_16),
    .ready_i_merge_pe               (merge_ready_i_8_16),

    .valid_i_gather_pe              (gather_valid_i_8_16),
    .data_i_gather_pe               (gather_data_i_8_16),
    .ready_o_gather_pe              (gather_ready_o_8_16),
    .valid_o_gather_pe              (gather_valid_o_8_16),
    .data_o_gather_pe               (gather_data_o_8_16),
    .ready_i_gather_pe              (gather_ready_i_8_16),

    .credit_upd                     (credit_upd[8][16])
);


network_interface #(
    .cast_out                       (cast_out_8_17),
    .gather_out                     (gather_out_8_17),
    .cast_sid                       (cast_sid_8_17),
    .gather_sid                     (gather_sid_8_17)
)ni_8_17(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[8][17]),
    .data_i_cast_nw                 (data_o_cast_nw[8][17]),
    .ready_o_cast_nw                (ready_i_cast_nw[8][17]),
    .valid_o_cast_nw                (valid_i_cast_nw[8][17]),
    .data_o_cast_nw                 (data_i_cast_nw[8][17]),
    .ready_i_cast_nw                (ready_o_cast_nw[8][17]),

    .valid_i_gather_nw              (valid_o_gather_nw[8][17]),
    .data_i_gather_nw               (data_o_gather_nw[8][17]),
    .ready_o_gather_nw              (ready_i_gather_nw[8][17]),
    .valid_o_gather_nw              (valid_i_gather_nw[8][17]),
    .data_o_gather_nw               (data_i_gather_nw[8][17]),
    .ready_i_gather_nw              (ready_o_gather_nw[8][17]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[8][17]),
    .data_i_merge_nw                (data_o_merge_nw[8][17]),
    .ready_o_merge_nw               (ready_i_merge_nw[8][17]),
    .valid_o_merge_nw               (valid_i_merge_nw[8][17]),
    .data_o_merge_nw                (data_i_merge_nw[8][17]),
    .ready_i_merge_nw               (ready_o_merge_nw[8][17]),

    .valid_i_cast_pe                (cast_valid_i_8_17),
    .data_i_cast_pe                 (cast_data_i_8_17),
    .ready_o_cast_pe                (cast_ready_o_8_17),
    .valid_o_cast_pe                (cast_valid_o_8_17),
    .data_o_cast_pe                 (cast_data_o_8_17),
    .ready_i_cast_pe                (cast_ready_i_8_17),

    .valid_i_merge_pe               (merge_valid_i_8_17),
    .data_i_merge_pe                (merge_data_i_8_17),
    .ready_o_merge_pe               (merge_ready_o_8_17),
    .valid_o_merge_pe               (merge_valid_o_8_17),
    .data_o_merge_pe                (merge_data_o_8_17),
    .ready_i_merge_pe               (merge_ready_i_8_17),

    .valid_i_gather_pe              (gather_valid_i_8_17),
    .data_i_gather_pe               (gather_data_i_8_17),
    .ready_o_gather_pe              (gather_ready_o_8_17),
    .valid_o_gather_pe              (gather_valid_o_8_17),
    .data_o_gather_pe               (gather_data_o_8_17),
    .ready_i_gather_pe              (gather_ready_i_8_17),

    .credit_upd                     (credit_upd[8][17])
);


network_interface #(
    .cast_out                       (cast_out_8_18),
    .gather_out                     (gather_out_8_18),
    .cast_sid                       (cast_sid_8_18),
    .gather_sid                     (gather_sid_8_18)
)ni_8_18(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[8][18]),
    .data_i_cast_nw                 (data_o_cast_nw[8][18]),
    .ready_o_cast_nw                (ready_i_cast_nw[8][18]),
    .valid_o_cast_nw                (valid_i_cast_nw[8][18]),
    .data_o_cast_nw                 (data_i_cast_nw[8][18]),
    .ready_i_cast_nw                (ready_o_cast_nw[8][18]),

    .valid_i_gather_nw              (valid_o_gather_nw[8][18]),
    .data_i_gather_nw               (data_o_gather_nw[8][18]),
    .ready_o_gather_nw              (ready_i_gather_nw[8][18]),
    .valid_o_gather_nw              (valid_i_gather_nw[8][18]),
    .data_o_gather_nw               (data_i_gather_nw[8][18]),
    .ready_i_gather_nw              (ready_o_gather_nw[8][18]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[8][18]),
    .data_i_merge_nw                (data_o_merge_nw[8][18]),
    .ready_o_merge_nw               (ready_i_merge_nw[8][18]),
    .valid_o_merge_nw               (valid_i_merge_nw[8][18]),
    .data_o_merge_nw                (data_i_merge_nw[8][18]),
    .ready_i_merge_nw               (ready_o_merge_nw[8][18]),

    .valid_i_cast_pe                (cast_valid_i_8_18),
    .data_i_cast_pe                 (cast_data_i_8_18),
    .ready_o_cast_pe                (cast_ready_o_8_18),
    .valid_o_cast_pe                (cast_valid_o_8_18),
    .data_o_cast_pe                 (cast_data_o_8_18),
    .ready_i_cast_pe                (cast_ready_i_8_18),

    .valid_i_merge_pe               (merge_valid_i_8_18),
    .data_i_merge_pe                (merge_data_i_8_18),
    .ready_o_merge_pe               (merge_ready_o_8_18),
    .valid_o_merge_pe               (merge_valid_o_8_18),
    .data_o_merge_pe                (merge_data_o_8_18),
    .ready_i_merge_pe               (merge_ready_i_8_18),

    .valid_i_gather_pe              (gather_valid_i_8_18),
    .data_i_gather_pe               (gather_data_i_8_18),
    .ready_o_gather_pe              (gather_ready_o_8_18),
    .valid_o_gather_pe              (gather_valid_o_8_18),
    .data_o_gather_pe               (gather_data_o_8_18),
    .ready_i_gather_pe              (gather_ready_i_8_18),

    .credit_upd                     (credit_upd[8][18])
);


network_interface #(
    .cast_out                       (cast_out_8_19),
    .gather_out                     (gather_out_8_19),
    .cast_sid                       (cast_sid_8_19),
    .gather_sid                     (gather_sid_8_19)
)ni_8_19(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[8][19]),
    .data_i_cast_nw                 (data_o_cast_nw[8][19]),
    .ready_o_cast_nw                (ready_i_cast_nw[8][19]),
    .valid_o_cast_nw                (valid_i_cast_nw[8][19]),
    .data_o_cast_nw                 (data_i_cast_nw[8][19]),
    .ready_i_cast_nw                (ready_o_cast_nw[8][19]),

    .valid_i_gather_nw              (valid_o_gather_nw[8][19]),
    .data_i_gather_nw               (data_o_gather_nw[8][19]),
    .ready_o_gather_nw              (ready_i_gather_nw[8][19]),
    .valid_o_gather_nw              (valid_i_gather_nw[8][19]),
    .data_o_gather_nw               (data_i_gather_nw[8][19]),
    .ready_i_gather_nw              (ready_o_gather_nw[8][19]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[8][19]),
    .data_i_merge_nw                (data_o_merge_nw[8][19]),
    .ready_o_merge_nw               (ready_i_merge_nw[8][19]),
    .valid_o_merge_nw               (valid_i_merge_nw[8][19]),
    .data_o_merge_nw                (data_i_merge_nw[8][19]),
    .ready_i_merge_nw               (ready_o_merge_nw[8][19]),

    .valid_i_cast_pe                (cast_valid_i_8_19),
    .data_i_cast_pe                 (cast_data_i_8_19),
    .ready_o_cast_pe                (cast_ready_o_8_19),
    .valid_o_cast_pe                (cast_valid_o_8_19),
    .data_o_cast_pe                 (cast_data_o_8_19),
    .ready_i_cast_pe                (cast_ready_i_8_19),

    .valid_i_merge_pe               (merge_valid_i_8_19),
    .data_i_merge_pe                (merge_data_i_8_19),
    .ready_o_merge_pe               (merge_ready_o_8_19),
    .valid_o_merge_pe               (merge_valid_o_8_19),
    .data_o_merge_pe                (merge_data_o_8_19),
    .ready_i_merge_pe               (merge_ready_i_8_19),

    .valid_i_gather_pe              (gather_valid_i_8_19),
    .data_i_gather_pe               (gather_data_i_8_19),
    .ready_o_gather_pe              (gather_ready_o_8_19),
    .valid_o_gather_pe              (gather_valid_o_8_19),
    .data_o_gather_pe               (gather_data_o_8_19),
    .ready_i_gather_pe              (gather_ready_i_8_19),

    .credit_upd                     (credit_upd[8][19])
);


network_interface #(
    .cast_out                       (cast_out_8_20),
    .gather_out                     (gather_out_8_20),
    .cast_sid                       (cast_sid_8_20),
    .gather_sid                     (gather_sid_8_20)
)ni_8_20(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[8][20]),
    .data_i_cast_nw                 (data_o_cast_nw[8][20]),
    .ready_o_cast_nw                (ready_i_cast_nw[8][20]),
    .valid_o_cast_nw                (valid_i_cast_nw[8][20]),
    .data_o_cast_nw                 (data_i_cast_nw[8][20]),
    .ready_i_cast_nw                (ready_o_cast_nw[8][20]),

    .valid_i_gather_nw              (valid_o_gather_nw[8][20]),
    .data_i_gather_nw               (data_o_gather_nw[8][20]),
    .ready_o_gather_nw              (ready_i_gather_nw[8][20]),
    .valid_o_gather_nw              (valid_i_gather_nw[8][20]),
    .data_o_gather_nw               (data_i_gather_nw[8][20]),
    .ready_i_gather_nw              (ready_o_gather_nw[8][20]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[8][20]),
    .data_i_merge_nw                (data_o_merge_nw[8][20]),
    .ready_o_merge_nw               (ready_i_merge_nw[8][20]),
    .valid_o_merge_nw               (valid_i_merge_nw[8][20]),
    .data_o_merge_nw                (data_i_merge_nw[8][20]),
    .ready_i_merge_nw               (ready_o_merge_nw[8][20]),

    .valid_i_cast_pe                (cast_valid_i_8_20),
    .data_i_cast_pe                 (cast_data_i_8_20),
    .ready_o_cast_pe                (cast_ready_o_8_20),
    .valid_o_cast_pe                (cast_valid_o_8_20),
    .data_o_cast_pe                 (cast_data_o_8_20),
    .ready_i_cast_pe                (cast_ready_i_8_20),

    .valid_i_merge_pe               (merge_valid_i_8_20),
    .data_i_merge_pe                (merge_data_i_8_20),
    .ready_o_merge_pe               (merge_ready_o_8_20),
    .valid_o_merge_pe               (merge_valid_o_8_20),
    .data_o_merge_pe                (merge_data_o_8_20),
    .ready_i_merge_pe               (merge_ready_i_8_20),

    .valid_i_gather_pe              (gather_valid_i_8_20),
    .data_i_gather_pe               (gather_data_i_8_20),
    .ready_o_gather_pe              (gather_ready_o_8_20),
    .valid_o_gather_pe              (gather_valid_o_8_20),
    .data_o_gather_pe               (gather_data_o_8_20),
    .ready_i_gather_pe              (gather_ready_i_8_20),

    .credit_upd                     (credit_upd[8][20])
);


network_interface #(
    .cast_out                       (cast_out_8_21),
    .gather_out                     (gather_out_8_21),
    .cast_sid                       (cast_sid_8_21),
    .gather_sid                     (gather_sid_8_21)
)ni_8_21(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[8][21]),
    .data_i_cast_nw                 (data_o_cast_nw[8][21]),
    .ready_o_cast_nw                (ready_i_cast_nw[8][21]),
    .valid_o_cast_nw                (valid_i_cast_nw[8][21]),
    .data_o_cast_nw                 (data_i_cast_nw[8][21]),
    .ready_i_cast_nw                (ready_o_cast_nw[8][21]),

    .valid_i_gather_nw              (valid_o_gather_nw[8][21]),
    .data_i_gather_nw               (data_o_gather_nw[8][21]),
    .ready_o_gather_nw              (ready_i_gather_nw[8][21]),
    .valid_o_gather_nw              (valid_i_gather_nw[8][21]),
    .data_o_gather_nw               (data_i_gather_nw[8][21]),
    .ready_i_gather_nw              (ready_o_gather_nw[8][21]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[8][21]),
    .data_i_merge_nw                (data_o_merge_nw[8][21]),
    .ready_o_merge_nw               (ready_i_merge_nw[8][21]),
    .valid_o_merge_nw               (valid_i_merge_nw[8][21]),
    .data_o_merge_nw                (data_i_merge_nw[8][21]),
    .ready_i_merge_nw               (ready_o_merge_nw[8][21]),

    .valid_i_cast_pe                (cast_valid_i_8_21),
    .data_i_cast_pe                 (cast_data_i_8_21),
    .ready_o_cast_pe                (cast_ready_o_8_21),
    .valid_o_cast_pe                (cast_valid_o_8_21),
    .data_o_cast_pe                 (cast_data_o_8_21),
    .ready_i_cast_pe                (cast_ready_i_8_21),

    .valid_i_merge_pe               (merge_valid_i_8_21),
    .data_i_merge_pe                (merge_data_i_8_21),
    .ready_o_merge_pe               (merge_ready_o_8_21),
    .valid_o_merge_pe               (merge_valid_o_8_21),
    .data_o_merge_pe                (merge_data_o_8_21),
    .ready_i_merge_pe               (merge_ready_i_8_21),

    .valid_i_gather_pe              (gather_valid_i_8_21),
    .data_i_gather_pe               (gather_data_i_8_21),
    .ready_o_gather_pe              (gather_ready_o_8_21),
    .valid_o_gather_pe              (gather_valid_o_8_21),
    .data_o_gather_pe               (gather_data_o_8_21),
    .ready_i_gather_pe              (gather_ready_i_8_21),

    .credit_upd                     (credit_upd[8][21])
);


network_interface #(
    .cast_out                       (cast_out_8_22),
    .gather_out                     (gather_out_8_22),
    .cast_sid                       (cast_sid_8_22),
    .gather_sid                     (gather_sid_8_22)
)ni_8_22(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[8][22]),
    .data_i_cast_nw                 (data_o_cast_nw[8][22]),
    .ready_o_cast_nw                (ready_i_cast_nw[8][22]),
    .valid_o_cast_nw                (valid_i_cast_nw[8][22]),
    .data_o_cast_nw                 (data_i_cast_nw[8][22]),
    .ready_i_cast_nw                (ready_o_cast_nw[8][22]),

    .valid_i_gather_nw              (valid_o_gather_nw[8][22]),
    .data_i_gather_nw               (data_o_gather_nw[8][22]),
    .ready_o_gather_nw              (ready_i_gather_nw[8][22]),
    .valid_o_gather_nw              (valid_i_gather_nw[8][22]),
    .data_o_gather_nw               (data_i_gather_nw[8][22]),
    .ready_i_gather_nw              (ready_o_gather_nw[8][22]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[8][22]),
    .data_i_merge_nw                (data_o_merge_nw[8][22]),
    .ready_o_merge_nw               (ready_i_merge_nw[8][22]),
    .valid_o_merge_nw               (valid_i_merge_nw[8][22]),
    .data_o_merge_nw                (data_i_merge_nw[8][22]),
    .ready_i_merge_nw               (ready_o_merge_nw[8][22]),

    .valid_i_cast_pe                (cast_valid_i_8_22),
    .data_i_cast_pe                 (cast_data_i_8_22),
    .ready_o_cast_pe                (cast_ready_o_8_22),
    .valid_o_cast_pe                (cast_valid_o_8_22),
    .data_o_cast_pe                 (cast_data_o_8_22),
    .ready_i_cast_pe                (cast_ready_i_8_22),

    .valid_i_merge_pe               (merge_valid_i_8_22),
    .data_i_merge_pe                (merge_data_i_8_22),
    .ready_o_merge_pe               (merge_ready_o_8_22),
    .valid_o_merge_pe               (merge_valid_o_8_22),
    .data_o_merge_pe                (merge_data_o_8_22),
    .ready_i_merge_pe               (merge_ready_i_8_22),

    .valid_i_gather_pe              (gather_valid_i_8_22),
    .data_i_gather_pe               (gather_data_i_8_22),
    .ready_o_gather_pe              (gather_ready_o_8_22),
    .valid_o_gather_pe              (gather_valid_o_8_22),
    .data_o_gather_pe               (gather_data_o_8_22),
    .ready_i_gather_pe              (gather_ready_i_8_22),

    .credit_upd                     (credit_upd[8][22])
);


network_interface #(
    .cast_out                       (cast_out_8_23),
    .gather_out                     (gather_out_8_23),
    .cast_sid                       (cast_sid_8_23),
    .gather_sid                     (gather_sid_8_23)
)ni_8_23(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[8][23]),
    .data_i_cast_nw                 (data_o_cast_nw[8][23]),
    .ready_o_cast_nw                (ready_i_cast_nw[8][23]),
    .valid_o_cast_nw                (valid_i_cast_nw[8][23]),
    .data_o_cast_nw                 (data_i_cast_nw[8][23]),
    .ready_i_cast_nw                (ready_o_cast_nw[8][23]),

    .valid_i_gather_nw              (valid_o_gather_nw[8][23]),
    .data_i_gather_nw               (data_o_gather_nw[8][23]),
    .ready_o_gather_nw              (ready_i_gather_nw[8][23]),
    .valid_o_gather_nw              (valid_i_gather_nw[8][23]),
    .data_o_gather_nw               (data_i_gather_nw[8][23]),
    .ready_i_gather_nw              (ready_o_gather_nw[8][23]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[8][23]),
    .data_i_merge_nw                (data_o_merge_nw[8][23]),
    .ready_o_merge_nw               (ready_i_merge_nw[8][23]),
    .valid_o_merge_nw               (valid_i_merge_nw[8][23]),
    .data_o_merge_nw                (data_i_merge_nw[8][23]),
    .ready_i_merge_nw               (ready_o_merge_nw[8][23]),

    .valid_i_cast_pe                (cast_valid_i_8_23),
    .data_i_cast_pe                 (cast_data_i_8_23),
    .ready_o_cast_pe                (cast_ready_o_8_23),
    .valid_o_cast_pe                (cast_valid_o_8_23),
    .data_o_cast_pe                 (cast_data_o_8_23),
    .ready_i_cast_pe                (cast_ready_i_8_23),

    .valid_i_merge_pe               (merge_valid_i_8_23),
    .data_i_merge_pe                (merge_data_i_8_23),
    .ready_o_merge_pe               (merge_ready_o_8_23),
    .valid_o_merge_pe               (merge_valid_o_8_23),
    .data_o_merge_pe                (merge_data_o_8_23),
    .ready_i_merge_pe               (merge_ready_i_8_23),

    .valid_i_gather_pe              (gather_valid_i_8_23),
    .data_i_gather_pe               (gather_data_i_8_23),
    .ready_o_gather_pe              (gather_ready_o_8_23),
    .valid_o_gather_pe              (gather_valid_o_8_23),
    .data_o_gather_pe               (gather_data_o_8_23),
    .ready_i_gather_pe              (gather_ready_i_8_23),

    .credit_upd                     (credit_upd[8][23])
);


network_interface #(
    .cast_out                       (cast_out_8_24),
    .gather_out                     (gather_out_8_24),
    .cast_sid                       (cast_sid_8_24),
    .gather_sid                     (gather_sid_8_24)
)ni_8_24(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[8][24]),
    .data_i_cast_nw                 (data_o_cast_nw[8][24]),
    .ready_o_cast_nw                (ready_i_cast_nw[8][24]),
    .valid_o_cast_nw                (valid_i_cast_nw[8][24]),
    .data_o_cast_nw                 (data_i_cast_nw[8][24]),
    .ready_i_cast_nw                (ready_o_cast_nw[8][24]),

    .valid_i_gather_nw              (valid_o_gather_nw[8][24]),
    .data_i_gather_nw               (data_o_gather_nw[8][24]),
    .ready_o_gather_nw              (ready_i_gather_nw[8][24]),
    .valid_o_gather_nw              (valid_i_gather_nw[8][24]),
    .data_o_gather_nw               (data_i_gather_nw[8][24]),
    .ready_i_gather_nw              (ready_o_gather_nw[8][24]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[8][24]),
    .data_i_merge_nw                (data_o_merge_nw[8][24]),
    .ready_o_merge_nw               (ready_i_merge_nw[8][24]),
    .valid_o_merge_nw               (valid_i_merge_nw[8][24]),
    .data_o_merge_nw                (data_i_merge_nw[8][24]),
    .ready_i_merge_nw               (ready_o_merge_nw[8][24]),

    .valid_i_cast_pe                (cast_valid_i_8_24),
    .data_i_cast_pe                 (cast_data_i_8_24),
    .ready_o_cast_pe                (cast_ready_o_8_24),
    .valid_o_cast_pe                (cast_valid_o_8_24),
    .data_o_cast_pe                 (cast_data_o_8_24),
    .ready_i_cast_pe                (cast_ready_i_8_24),

    .valid_i_merge_pe               (merge_valid_i_8_24),
    .data_i_merge_pe                (merge_data_i_8_24),
    .ready_o_merge_pe               (merge_ready_o_8_24),
    .valid_o_merge_pe               (merge_valid_o_8_24),
    .data_o_merge_pe                (merge_data_o_8_24),
    .ready_i_merge_pe               (merge_ready_i_8_24),

    .valid_i_gather_pe              (gather_valid_i_8_24),
    .data_i_gather_pe               (gather_data_i_8_24),
    .ready_o_gather_pe              (gather_ready_o_8_24),
    .valid_o_gather_pe              (gather_valid_o_8_24),
    .data_o_gather_pe               (gather_data_o_8_24),
    .ready_i_gather_pe              (gather_ready_i_8_24),

    .credit_upd                     (credit_upd[8][24])
);


network_interface #(
    .cast_out                       (cast_out_9_0),
    .gather_out                     (gather_out_9_0),
    .cast_sid                       (cast_sid_9_0),
    .gather_sid                     (gather_sid_9_0)
)ni_9_0(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[9][0]),
    .data_i_cast_nw                 (data_o_cast_nw[9][0]),
    .ready_o_cast_nw                (ready_i_cast_nw[9][0]),
    .valid_o_cast_nw                (valid_i_cast_nw[9][0]),
    .data_o_cast_nw                 (data_i_cast_nw[9][0]),
    .ready_i_cast_nw                (ready_o_cast_nw[9][0]),

    .valid_i_gather_nw              (valid_o_gather_nw[9][0]),
    .data_i_gather_nw               (data_o_gather_nw[9][0]),
    .ready_o_gather_nw              (ready_i_gather_nw[9][0]),
    .valid_o_gather_nw              (valid_i_gather_nw[9][0]),
    .data_o_gather_nw               (data_i_gather_nw[9][0]),
    .ready_i_gather_nw              (ready_o_gather_nw[9][0]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[9][0]),
    .data_i_merge_nw                (data_o_merge_nw[9][0]),
    .ready_o_merge_nw               (ready_i_merge_nw[9][0]),
    .valid_o_merge_nw               (valid_i_merge_nw[9][0]),
    .data_o_merge_nw                (data_i_merge_nw[9][0]),
    .ready_i_merge_nw               (ready_o_merge_nw[9][0]),

    .valid_i_cast_pe                (cast_valid_i_9_0),
    .data_i_cast_pe                 (cast_data_i_9_0),
    .ready_o_cast_pe                (cast_ready_o_9_0),
    .valid_o_cast_pe                (cast_valid_o_9_0),
    .data_o_cast_pe                 (cast_data_o_9_0),
    .ready_i_cast_pe                (cast_ready_i_9_0),

    .valid_i_merge_pe               (merge_valid_i_9_0),
    .data_i_merge_pe                (merge_data_i_9_0),
    .ready_o_merge_pe               (merge_ready_o_9_0),
    .valid_o_merge_pe               (merge_valid_o_9_0),
    .data_o_merge_pe                (merge_data_o_9_0),
    .ready_i_merge_pe               (merge_ready_i_9_0),

    .valid_i_gather_pe              (gather_valid_i_9_0),
    .data_i_gather_pe               (gather_data_i_9_0),
    .ready_o_gather_pe              (gather_ready_o_9_0),
    .valid_o_gather_pe              (gather_valid_o_9_0),
    .data_o_gather_pe               (gather_data_o_9_0),
    .ready_i_gather_pe              (gather_ready_i_9_0),

    .credit_upd                     (credit_upd[9][0])
);


network_interface #(
    .cast_out                       (cast_out_9_1),
    .gather_out                     (gather_out_9_1),
    .cast_sid                       (cast_sid_9_1),
    .gather_sid                     (gather_sid_9_1)
)ni_9_1(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[9][1]),
    .data_i_cast_nw                 (data_o_cast_nw[9][1]),
    .ready_o_cast_nw                (ready_i_cast_nw[9][1]),
    .valid_o_cast_nw                (valid_i_cast_nw[9][1]),
    .data_o_cast_nw                 (data_i_cast_nw[9][1]),
    .ready_i_cast_nw                (ready_o_cast_nw[9][1]),

    .valid_i_gather_nw              (valid_o_gather_nw[9][1]),
    .data_i_gather_nw               (data_o_gather_nw[9][1]),
    .ready_o_gather_nw              (ready_i_gather_nw[9][1]),
    .valid_o_gather_nw              (valid_i_gather_nw[9][1]),
    .data_o_gather_nw               (data_i_gather_nw[9][1]),
    .ready_i_gather_nw              (ready_o_gather_nw[9][1]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[9][1]),
    .data_i_merge_nw                (data_o_merge_nw[9][1]),
    .ready_o_merge_nw               (ready_i_merge_nw[9][1]),
    .valid_o_merge_nw               (valid_i_merge_nw[9][1]),
    .data_o_merge_nw                (data_i_merge_nw[9][1]),
    .ready_i_merge_nw               (ready_o_merge_nw[9][1]),

    .valid_i_cast_pe                (cast_valid_i_9_1),
    .data_i_cast_pe                 (cast_data_i_9_1),
    .ready_o_cast_pe                (cast_ready_o_9_1),
    .valid_o_cast_pe                (cast_valid_o_9_1),
    .data_o_cast_pe                 (cast_data_o_9_1),
    .ready_i_cast_pe                (cast_ready_i_9_1),

    .valid_i_merge_pe               (merge_valid_i_9_1),
    .data_i_merge_pe                (merge_data_i_9_1),
    .ready_o_merge_pe               (merge_ready_o_9_1),
    .valid_o_merge_pe               (merge_valid_o_9_1),
    .data_o_merge_pe                (merge_data_o_9_1),
    .ready_i_merge_pe               (merge_ready_i_9_1),

    .valid_i_gather_pe              (gather_valid_i_9_1),
    .data_i_gather_pe               (gather_data_i_9_1),
    .ready_o_gather_pe              (gather_ready_o_9_1),
    .valid_o_gather_pe              (gather_valid_o_9_1),
    .data_o_gather_pe               (gather_data_o_9_1),
    .ready_i_gather_pe              (gather_ready_i_9_1),

    .credit_upd                     (credit_upd[9][1])
);


network_interface #(
    .cast_out                       (cast_out_9_2),
    .gather_out                     (gather_out_9_2),
    .cast_sid                       (cast_sid_9_2),
    .gather_sid                     (gather_sid_9_2)
)ni_9_2(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[9][2]),
    .data_i_cast_nw                 (data_o_cast_nw[9][2]),
    .ready_o_cast_nw                (ready_i_cast_nw[9][2]),
    .valid_o_cast_nw                (valid_i_cast_nw[9][2]),
    .data_o_cast_nw                 (data_i_cast_nw[9][2]),
    .ready_i_cast_nw                (ready_o_cast_nw[9][2]),

    .valid_i_gather_nw              (valid_o_gather_nw[9][2]),
    .data_i_gather_nw               (data_o_gather_nw[9][2]),
    .ready_o_gather_nw              (ready_i_gather_nw[9][2]),
    .valid_o_gather_nw              (valid_i_gather_nw[9][2]),
    .data_o_gather_nw               (data_i_gather_nw[9][2]),
    .ready_i_gather_nw              (ready_o_gather_nw[9][2]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[9][2]),
    .data_i_merge_nw                (data_o_merge_nw[9][2]),
    .ready_o_merge_nw               (ready_i_merge_nw[9][2]),
    .valid_o_merge_nw               (valid_i_merge_nw[9][2]),
    .data_o_merge_nw                (data_i_merge_nw[9][2]),
    .ready_i_merge_nw               (ready_o_merge_nw[9][2]),

    .valid_i_cast_pe                (cast_valid_i_9_2),
    .data_i_cast_pe                 (cast_data_i_9_2),
    .ready_o_cast_pe                (cast_ready_o_9_2),
    .valid_o_cast_pe                (cast_valid_o_9_2),
    .data_o_cast_pe                 (cast_data_o_9_2),
    .ready_i_cast_pe                (cast_ready_i_9_2),

    .valid_i_merge_pe               (merge_valid_i_9_2),
    .data_i_merge_pe                (merge_data_i_9_2),
    .ready_o_merge_pe               (merge_ready_o_9_2),
    .valid_o_merge_pe               (merge_valid_o_9_2),
    .data_o_merge_pe                (merge_data_o_9_2),
    .ready_i_merge_pe               (merge_ready_i_9_2),

    .valid_i_gather_pe              (gather_valid_i_9_2),
    .data_i_gather_pe               (gather_data_i_9_2),
    .ready_o_gather_pe              (gather_ready_o_9_2),
    .valid_o_gather_pe              (gather_valid_o_9_2),
    .data_o_gather_pe               (gather_data_o_9_2),
    .ready_i_gather_pe              (gather_ready_i_9_2),

    .credit_upd                     (credit_upd[9][2])
);


network_interface #(
    .cast_out                       (cast_out_9_3),
    .gather_out                     (gather_out_9_3),
    .cast_sid                       (cast_sid_9_3),
    .gather_sid                     (gather_sid_9_3)
)ni_9_3(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[9][3]),
    .data_i_cast_nw                 (data_o_cast_nw[9][3]),
    .ready_o_cast_nw                (ready_i_cast_nw[9][3]),
    .valid_o_cast_nw                (valid_i_cast_nw[9][3]),
    .data_o_cast_nw                 (data_i_cast_nw[9][3]),
    .ready_i_cast_nw                (ready_o_cast_nw[9][3]),

    .valid_i_gather_nw              (valid_o_gather_nw[9][3]),
    .data_i_gather_nw               (data_o_gather_nw[9][3]),
    .ready_o_gather_nw              (ready_i_gather_nw[9][3]),
    .valid_o_gather_nw              (valid_i_gather_nw[9][3]),
    .data_o_gather_nw               (data_i_gather_nw[9][3]),
    .ready_i_gather_nw              (ready_o_gather_nw[9][3]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[9][3]),
    .data_i_merge_nw                (data_o_merge_nw[9][3]),
    .ready_o_merge_nw               (ready_i_merge_nw[9][3]),
    .valid_o_merge_nw               (valid_i_merge_nw[9][3]),
    .data_o_merge_nw                (data_i_merge_nw[9][3]),
    .ready_i_merge_nw               (ready_o_merge_nw[9][3]),

    .valid_i_cast_pe                (cast_valid_i_9_3),
    .data_i_cast_pe                 (cast_data_i_9_3),
    .ready_o_cast_pe                (cast_ready_o_9_3),
    .valid_o_cast_pe                (cast_valid_o_9_3),
    .data_o_cast_pe                 (cast_data_o_9_3),
    .ready_i_cast_pe                (cast_ready_i_9_3),

    .valid_i_merge_pe               (merge_valid_i_9_3),
    .data_i_merge_pe                (merge_data_i_9_3),
    .ready_o_merge_pe               (merge_ready_o_9_3),
    .valid_o_merge_pe               (merge_valid_o_9_3),
    .data_o_merge_pe                (merge_data_o_9_3),
    .ready_i_merge_pe               (merge_ready_i_9_3),

    .valid_i_gather_pe              (gather_valid_i_9_3),
    .data_i_gather_pe               (gather_data_i_9_3),
    .ready_o_gather_pe              (gather_ready_o_9_3),
    .valid_o_gather_pe              (gather_valid_o_9_3),
    .data_o_gather_pe               (gather_data_o_9_3),
    .ready_i_gather_pe              (gather_ready_i_9_3),

    .credit_upd                     (credit_upd[9][3])
);


network_interface #(
    .cast_out                       (cast_out_9_4),
    .gather_out                     (gather_out_9_4),
    .cast_sid                       (cast_sid_9_4),
    .gather_sid                     (gather_sid_9_4)
)ni_9_4(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[9][4]),
    .data_i_cast_nw                 (data_o_cast_nw[9][4]),
    .ready_o_cast_nw                (ready_i_cast_nw[9][4]),
    .valid_o_cast_nw                (valid_i_cast_nw[9][4]),
    .data_o_cast_nw                 (data_i_cast_nw[9][4]),
    .ready_i_cast_nw                (ready_o_cast_nw[9][4]),

    .valid_i_gather_nw              (valid_o_gather_nw[9][4]),
    .data_i_gather_nw               (data_o_gather_nw[9][4]),
    .ready_o_gather_nw              (ready_i_gather_nw[9][4]),
    .valid_o_gather_nw              (valid_i_gather_nw[9][4]),
    .data_o_gather_nw               (data_i_gather_nw[9][4]),
    .ready_i_gather_nw              (ready_o_gather_nw[9][4]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[9][4]),
    .data_i_merge_nw                (data_o_merge_nw[9][4]),
    .ready_o_merge_nw               (ready_i_merge_nw[9][4]),
    .valid_o_merge_nw               (valid_i_merge_nw[9][4]),
    .data_o_merge_nw                (data_i_merge_nw[9][4]),
    .ready_i_merge_nw               (ready_o_merge_nw[9][4]),

    .valid_i_cast_pe                (cast_valid_i_9_4),
    .data_i_cast_pe                 (cast_data_i_9_4),
    .ready_o_cast_pe                (cast_ready_o_9_4),
    .valid_o_cast_pe                (cast_valid_o_9_4),
    .data_o_cast_pe                 (cast_data_o_9_4),
    .ready_i_cast_pe                (cast_ready_i_9_4),

    .valid_i_merge_pe               (merge_valid_i_9_4),
    .data_i_merge_pe                (merge_data_i_9_4),
    .ready_o_merge_pe               (merge_ready_o_9_4),
    .valid_o_merge_pe               (merge_valid_o_9_4),
    .data_o_merge_pe                (merge_data_o_9_4),
    .ready_i_merge_pe               (merge_ready_i_9_4),

    .valid_i_gather_pe              (gather_valid_i_9_4),
    .data_i_gather_pe               (gather_data_i_9_4),
    .ready_o_gather_pe              (gather_ready_o_9_4),
    .valid_o_gather_pe              (gather_valid_o_9_4),
    .data_o_gather_pe               (gather_data_o_9_4),
    .ready_i_gather_pe              (gather_ready_i_9_4),

    .credit_upd                     (credit_upd[9][4])
);


network_interface #(
    .cast_out                       (cast_out_9_5),
    .gather_out                     (gather_out_9_5),
    .cast_sid                       (cast_sid_9_5),
    .gather_sid                     (gather_sid_9_5)
)ni_9_5(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[9][5]),
    .data_i_cast_nw                 (data_o_cast_nw[9][5]),
    .ready_o_cast_nw                (ready_i_cast_nw[9][5]),
    .valid_o_cast_nw                (valid_i_cast_nw[9][5]),
    .data_o_cast_nw                 (data_i_cast_nw[9][5]),
    .ready_i_cast_nw                (ready_o_cast_nw[9][5]),

    .valid_i_gather_nw              (valid_o_gather_nw[9][5]),
    .data_i_gather_nw               (data_o_gather_nw[9][5]),
    .ready_o_gather_nw              (ready_i_gather_nw[9][5]),
    .valid_o_gather_nw              (valid_i_gather_nw[9][5]),
    .data_o_gather_nw               (data_i_gather_nw[9][5]),
    .ready_i_gather_nw              (ready_o_gather_nw[9][5]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[9][5]),
    .data_i_merge_nw                (data_o_merge_nw[9][5]),
    .ready_o_merge_nw               (ready_i_merge_nw[9][5]),
    .valid_o_merge_nw               (valid_i_merge_nw[9][5]),
    .data_o_merge_nw                (data_i_merge_nw[9][5]),
    .ready_i_merge_nw               (ready_o_merge_nw[9][5]),

    .valid_i_cast_pe                (cast_valid_i_9_5),
    .data_i_cast_pe                 (cast_data_i_9_5),
    .ready_o_cast_pe                (cast_ready_o_9_5),
    .valid_o_cast_pe                (cast_valid_o_9_5),
    .data_o_cast_pe                 (cast_data_o_9_5),
    .ready_i_cast_pe                (cast_ready_i_9_5),

    .valid_i_merge_pe               (merge_valid_i_9_5),
    .data_i_merge_pe                (merge_data_i_9_5),
    .ready_o_merge_pe               (merge_ready_o_9_5),
    .valid_o_merge_pe               (merge_valid_o_9_5),
    .data_o_merge_pe                (merge_data_o_9_5),
    .ready_i_merge_pe               (merge_ready_i_9_5),

    .valid_i_gather_pe              (gather_valid_i_9_5),
    .data_i_gather_pe               (gather_data_i_9_5),
    .ready_o_gather_pe              (gather_ready_o_9_5),
    .valid_o_gather_pe              (gather_valid_o_9_5),
    .data_o_gather_pe               (gather_data_o_9_5),
    .ready_i_gather_pe              (gather_ready_i_9_5),

    .credit_upd                     (credit_upd[9][5])
);


network_interface #(
    .cast_out                       (cast_out_9_6),
    .gather_out                     (gather_out_9_6),
    .cast_sid                       (cast_sid_9_6),
    .gather_sid                     (gather_sid_9_6)
)ni_9_6(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[9][6]),
    .data_i_cast_nw                 (data_o_cast_nw[9][6]),
    .ready_o_cast_nw                (ready_i_cast_nw[9][6]),
    .valid_o_cast_nw                (valid_i_cast_nw[9][6]),
    .data_o_cast_nw                 (data_i_cast_nw[9][6]),
    .ready_i_cast_nw                (ready_o_cast_nw[9][6]),

    .valid_i_gather_nw              (valid_o_gather_nw[9][6]),
    .data_i_gather_nw               (data_o_gather_nw[9][6]),
    .ready_o_gather_nw              (ready_i_gather_nw[9][6]),
    .valid_o_gather_nw              (valid_i_gather_nw[9][6]),
    .data_o_gather_nw               (data_i_gather_nw[9][6]),
    .ready_i_gather_nw              (ready_o_gather_nw[9][6]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[9][6]),
    .data_i_merge_nw                (data_o_merge_nw[9][6]),
    .ready_o_merge_nw               (ready_i_merge_nw[9][6]),
    .valid_o_merge_nw               (valid_i_merge_nw[9][6]),
    .data_o_merge_nw                (data_i_merge_nw[9][6]),
    .ready_i_merge_nw               (ready_o_merge_nw[9][6]),

    .valid_i_cast_pe                (cast_valid_i_9_6),
    .data_i_cast_pe                 (cast_data_i_9_6),
    .ready_o_cast_pe                (cast_ready_o_9_6),
    .valid_o_cast_pe                (cast_valid_o_9_6),
    .data_o_cast_pe                 (cast_data_o_9_6),
    .ready_i_cast_pe                (cast_ready_i_9_6),

    .valid_i_merge_pe               (merge_valid_i_9_6),
    .data_i_merge_pe                (merge_data_i_9_6),
    .ready_o_merge_pe               (merge_ready_o_9_6),
    .valid_o_merge_pe               (merge_valid_o_9_6),
    .data_o_merge_pe                (merge_data_o_9_6),
    .ready_i_merge_pe               (merge_ready_i_9_6),

    .valid_i_gather_pe              (gather_valid_i_9_6),
    .data_i_gather_pe               (gather_data_i_9_6),
    .ready_o_gather_pe              (gather_ready_o_9_6),
    .valid_o_gather_pe              (gather_valid_o_9_6),
    .data_o_gather_pe               (gather_data_o_9_6),
    .ready_i_gather_pe              (gather_ready_i_9_6),

    .credit_upd                     (credit_upd[9][6])
);


network_interface #(
    .cast_out                       (cast_out_9_7),
    .gather_out                     (gather_out_9_7),
    .cast_sid                       (cast_sid_9_7),
    .gather_sid                     (gather_sid_9_7)
)ni_9_7(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[9][7]),
    .data_i_cast_nw                 (data_o_cast_nw[9][7]),
    .ready_o_cast_nw                (ready_i_cast_nw[9][7]),
    .valid_o_cast_nw                (valid_i_cast_nw[9][7]),
    .data_o_cast_nw                 (data_i_cast_nw[9][7]),
    .ready_i_cast_nw                (ready_o_cast_nw[9][7]),

    .valid_i_gather_nw              (valid_o_gather_nw[9][7]),
    .data_i_gather_nw               (data_o_gather_nw[9][7]),
    .ready_o_gather_nw              (ready_i_gather_nw[9][7]),
    .valid_o_gather_nw              (valid_i_gather_nw[9][7]),
    .data_o_gather_nw               (data_i_gather_nw[9][7]),
    .ready_i_gather_nw              (ready_o_gather_nw[9][7]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[9][7]),
    .data_i_merge_nw                (data_o_merge_nw[9][7]),
    .ready_o_merge_nw               (ready_i_merge_nw[9][7]),
    .valid_o_merge_nw               (valid_i_merge_nw[9][7]),
    .data_o_merge_nw                (data_i_merge_nw[9][7]),
    .ready_i_merge_nw               (ready_o_merge_nw[9][7]),

    .valid_i_cast_pe                (cast_valid_i_9_7),
    .data_i_cast_pe                 (cast_data_i_9_7),
    .ready_o_cast_pe                (cast_ready_o_9_7),
    .valid_o_cast_pe                (cast_valid_o_9_7),
    .data_o_cast_pe                 (cast_data_o_9_7),
    .ready_i_cast_pe                (cast_ready_i_9_7),

    .valid_i_merge_pe               (merge_valid_i_9_7),
    .data_i_merge_pe                (merge_data_i_9_7),
    .ready_o_merge_pe               (merge_ready_o_9_7),
    .valid_o_merge_pe               (merge_valid_o_9_7),
    .data_o_merge_pe                (merge_data_o_9_7),
    .ready_i_merge_pe               (merge_ready_i_9_7),

    .valid_i_gather_pe              (gather_valid_i_9_7),
    .data_i_gather_pe               (gather_data_i_9_7),
    .ready_o_gather_pe              (gather_ready_o_9_7),
    .valid_o_gather_pe              (gather_valid_o_9_7),
    .data_o_gather_pe               (gather_data_o_9_7),
    .ready_i_gather_pe              (gather_ready_i_9_7),

    .credit_upd                     (credit_upd[9][7])
);


network_interface #(
    .cast_out                       (cast_out_9_8),
    .gather_out                     (gather_out_9_8),
    .cast_sid                       (cast_sid_9_8),
    .gather_sid                     (gather_sid_9_8)
)ni_9_8(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[9][8]),
    .data_i_cast_nw                 (data_o_cast_nw[9][8]),
    .ready_o_cast_nw                (ready_i_cast_nw[9][8]),
    .valid_o_cast_nw                (valid_i_cast_nw[9][8]),
    .data_o_cast_nw                 (data_i_cast_nw[9][8]),
    .ready_i_cast_nw                (ready_o_cast_nw[9][8]),

    .valid_i_gather_nw              (valid_o_gather_nw[9][8]),
    .data_i_gather_nw               (data_o_gather_nw[9][8]),
    .ready_o_gather_nw              (ready_i_gather_nw[9][8]),
    .valid_o_gather_nw              (valid_i_gather_nw[9][8]),
    .data_o_gather_nw               (data_i_gather_nw[9][8]),
    .ready_i_gather_nw              (ready_o_gather_nw[9][8]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[9][8]),
    .data_i_merge_nw                (data_o_merge_nw[9][8]),
    .ready_o_merge_nw               (ready_i_merge_nw[9][8]),
    .valid_o_merge_nw               (valid_i_merge_nw[9][8]),
    .data_o_merge_nw                (data_i_merge_nw[9][8]),
    .ready_i_merge_nw               (ready_o_merge_nw[9][8]),

    .valid_i_cast_pe                (cast_valid_i_9_8),
    .data_i_cast_pe                 (cast_data_i_9_8),
    .ready_o_cast_pe                (cast_ready_o_9_8),
    .valid_o_cast_pe                (cast_valid_o_9_8),
    .data_o_cast_pe                 (cast_data_o_9_8),
    .ready_i_cast_pe                (cast_ready_i_9_8),

    .valid_i_merge_pe               (merge_valid_i_9_8),
    .data_i_merge_pe                (merge_data_i_9_8),
    .ready_o_merge_pe               (merge_ready_o_9_8),
    .valid_o_merge_pe               (merge_valid_o_9_8),
    .data_o_merge_pe                (merge_data_o_9_8),
    .ready_i_merge_pe               (merge_ready_i_9_8),

    .valid_i_gather_pe              (gather_valid_i_9_8),
    .data_i_gather_pe               (gather_data_i_9_8),
    .ready_o_gather_pe              (gather_ready_o_9_8),
    .valid_o_gather_pe              (gather_valid_o_9_8),
    .data_o_gather_pe               (gather_data_o_9_8),
    .ready_i_gather_pe              (gather_ready_i_9_8),

    .credit_upd                     (credit_upd[9][8])
);


network_interface #(
    .cast_out                       (cast_out_9_9),
    .gather_out                     (gather_out_9_9),
    .cast_sid                       (cast_sid_9_9),
    .gather_sid                     (gather_sid_9_9)
)ni_9_9(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[9][9]),
    .data_i_cast_nw                 (data_o_cast_nw[9][9]),
    .ready_o_cast_nw                (ready_i_cast_nw[9][9]),
    .valid_o_cast_nw                (valid_i_cast_nw[9][9]),
    .data_o_cast_nw                 (data_i_cast_nw[9][9]),
    .ready_i_cast_nw                (ready_o_cast_nw[9][9]),

    .valid_i_gather_nw              (valid_o_gather_nw[9][9]),
    .data_i_gather_nw               (data_o_gather_nw[9][9]),
    .ready_o_gather_nw              (ready_i_gather_nw[9][9]),
    .valid_o_gather_nw              (valid_i_gather_nw[9][9]),
    .data_o_gather_nw               (data_i_gather_nw[9][9]),
    .ready_i_gather_nw              (ready_o_gather_nw[9][9]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[9][9]),
    .data_i_merge_nw                (data_o_merge_nw[9][9]),
    .ready_o_merge_nw               (ready_i_merge_nw[9][9]),
    .valid_o_merge_nw               (valid_i_merge_nw[9][9]),
    .data_o_merge_nw                (data_i_merge_nw[9][9]),
    .ready_i_merge_nw               (ready_o_merge_nw[9][9]),

    .valid_i_cast_pe                (cast_valid_i_9_9),
    .data_i_cast_pe                 (cast_data_i_9_9),
    .ready_o_cast_pe                (cast_ready_o_9_9),
    .valid_o_cast_pe                (cast_valid_o_9_9),
    .data_o_cast_pe                 (cast_data_o_9_9),
    .ready_i_cast_pe                (cast_ready_i_9_9),

    .valid_i_merge_pe               (merge_valid_i_9_9),
    .data_i_merge_pe                (merge_data_i_9_9),
    .ready_o_merge_pe               (merge_ready_o_9_9),
    .valid_o_merge_pe               (merge_valid_o_9_9),
    .data_o_merge_pe                (merge_data_o_9_9),
    .ready_i_merge_pe               (merge_ready_i_9_9),

    .valid_i_gather_pe              (gather_valid_i_9_9),
    .data_i_gather_pe               (gather_data_i_9_9),
    .ready_o_gather_pe              (gather_ready_o_9_9),
    .valid_o_gather_pe              (gather_valid_o_9_9),
    .data_o_gather_pe               (gather_data_o_9_9),
    .ready_i_gather_pe              (gather_ready_i_9_9),

    .credit_upd                     (credit_upd[9][9])
);


network_interface #(
    .cast_out                       (cast_out_9_10),
    .gather_out                     (gather_out_9_10),
    .cast_sid                       (cast_sid_9_10),
    .gather_sid                     (gather_sid_9_10)
)ni_9_10(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[9][10]),
    .data_i_cast_nw                 (data_o_cast_nw[9][10]),
    .ready_o_cast_nw                (ready_i_cast_nw[9][10]),
    .valid_o_cast_nw                (valid_i_cast_nw[9][10]),
    .data_o_cast_nw                 (data_i_cast_nw[9][10]),
    .ready_i_cast_nw                (ready_o_cast_nw[9][10]),

    .valid_i_gather_nw              (valid_o_gather_nw[9][10]),
    .data_i_gather_nw               (data_o_gather_nw[9][10]),
    .ready_o_gather_nw              (ready_i_gather_nw[9][10]),
    .valid_o_gather_nw              (valid_i_gather_nw[9][10]),
    .data_o_gather_nw               (data_i_gather_nw[9][10]),
    .ready_i_gather_nw              (ready_o_gather_nw[9][10]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[9][10]),
    .data_i_merge_nw                (data_o_merge_nw[9][10]),
    .ready_o_merge_nw               (ready_i_merge_nw[9][10]),
    .valid_o_merge_nw               (valid_i_merge_nw[9][10]),
    .data_o_merge_nw                (data_i_merge_nw[9][10]),
    .ready_i_merge_nw               (ready_o_merge_nw[9][10]),

    .valid_i_cast_pe                (cast_valid_i_9_10),
    .data_i_cast_pe                 (cast_data_i_9_10),
    .ready_o_cast_pe                (cast_ready_o_9_10),
    .valid_o_cast_pe                (cast_valid_o_9_10),
    .data_o_cast_pe                 (cast_data_o_9_10),
    .ready_i_cast_pe                (cast_ready_i_9_10),

    .valid_i_merge_pe               (merge_valid_i_9_10),
    .data_i_merge_pe                (merge_data_i_9_10),
    .ready_o_merge_pe               (merge_ready_o_9_10),
    .valid_o_merge_pe               (merge_valid_o_9_10),
    .data_o_merge_pe                (merge_data_o_9_10),
    .ready_i_merge_pe               (merge_ready_i_9_10),

    .valid_i_gather_pe              (gather_valid_i_9_10),
    .data_i_gather_pe               (gather_data_i_9_10),
    .ready_o_gather_pe              (gather_ready_o_9_10),
    .valid_o_gather_pe              (gather_valid_o_9_10),
    .data_o_gather_pe               (gather_data_o_9_10),
    .ready_i_gather_pe              (gather_ready_i_9_10),

    .credit_upd                     (credit_upd[9][10])
);


network_interface #(
    .cast_out                       (cast_out_9_11),
    .gather_out                     (gather_out_9_11),
    .cast_sid                       (cast_sid_9_11),
    .gather_sid                     (gather_sid_9_11)
)ni_9_11(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[9][11]),
    .data_i_cast_nw                 (data_o_cast_nw[9][11]),
    .ready_o_cast_nw                (ready_i_cast_nw[9][11]),
    .valid_o_cast_nw                (valid_i_cast_nw[9][11]),
    .data_o_cast_nw                 (data_i_cast_nw[9][11]),
    .ready_i_cast_nw                (ready_o_cast_nw[9][11]),

    .valid_i_gather_nw              (valid_o_gather_nw[9][11]),
    .data_i_gather_nw               (data_o_gather_nw[9][11]),
    .ready_o_gather_nw              (ready_i_gather_nw[9][11]),
    .valid_o_gather_nw              (valid_i_gather_nw[9][11]),
    .data_o_gather_nw               (data_i_gather_nw[9][11]),
    .ready_i_gather_nw              (ready_o_gather_nw[9][11]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[9][11]),
    .data_i_merge_nw                (data_o_merge_nw[9][11]),
    .ready_o_merge_nw               (ready_i_merge_nw[9][11]),
    .valid_o_merge_nw               (valid_i_merge_nw[9][11]),
    .data_o_merge_nw                (data_i_merge_nw[9][11]),
    .ready_i_merge_nw               (ready_o_merge_nw[9][11]),

    .valid_i_cast_pe                (cast_valid_i_9_11),
    .data_i_cast_pe                 (cast_data_i_9_11),
    .ready_o_cast_pe                (cast_ready_o_9_11),
    .valid_o_cast_pe                (cast_valid_o_9_11),
    .data_o_cast_pe                 (cast_data_o_9_11),
    .ready_i_cast_pe                (cast_ready_i_9_11),

    .valid_i_merge_pe               (merge_valid_i_9_11),
    .data_i_merge_pe                (merge_data_i_9_11),
    .ready_o_merge_pe               (merge_ready_o_9_11),
    .valid_o_merge_pe               (merge_valid_o_9_11),
    .data_o_merge_pe                (merge_data_o_9_11),
    .ready_i_merge_pe               (merge_ready_i_9_11),

    .valid_i_gather_pe              (gather_valid_i_9_11),
    .data_i_gather_pe               (gather_data_i_9_11),
    .ready_o_gather_pe              (gather_ready_o_9_11),
    .valid_o_gather_pe              (gather_valid_o_9_11),
    .data_o_gather_pe               (gather_data_o_9_11),
    .ready_i_gather_pe              (gather_ready_i_9_11),

    .credit_upd                     (credit_upd[9][11])
);


network_interface #(
    .cast_out                       (cast_out_9_12),
    .gather_out                     (gather_out_9_12),
    .cast_sid                       (cast_sid_9_12),
    .gather_sid                     (gather_sid_9_12)
)ni_9_12(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[9][12]),
    .data_i_cast_nw                 (data_o_cast_nw[9][12]),
    .ready_o_cast_nw                (ready_i_cast_nw[9][12]),
    .valid_o_cast_nw                (valid_i_cast_nw[9][12]),
    .data_o_cast_nw                 (data_i_cast_nw[9][12]),
    .ready_i_cast_nw                (ready_o_cast_nw[9][12]),

    .valid_i_gather_nw              (valid_o_gather_nw[9][12]),
    .data_i_gather_nw               (data_o_gather_nw[9][12]),
    .ready_o_gather_nw              (ready_i_gather_nw[9][12]),
    .valid_o_gather_nw              (valid_i_gather_nw[9][12]),
    .data_o_gather_nw               (data_i_gather_nw[9][12]),
    .ready_i_gather_nw              (ready_o_gather_nw[9][12]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[9][12]),
    .data_i_merge_nw                (data_o_merge_nw[9][12]),
    .ready_o_merge_nw               (ready_i_merge_nw[9][12]),
    .valid_o_merge_nw               (valid_i_merge_nw[9][12]),
    .data_o_merge_nw                (data_i_merge_nw[9][12]),
    .ready_i_merge_nw               (ready_o_merge_nw[9][12]),

    .valid_i_cast_pe                (cast_valid_i_9_12),
    .data_i_cast_pe                 (cast_data_i_9_12),
    .ready_o_cast_pe                (cast_ready_o_9_12),
    .valid_o_cast_pe                (cast_valid_o_9_12),
    .data_o_cast_pe                 (cast_data_o_9_12),
    .ready_i_cast_pe                (cast_ready_i_9_12),

    .valid_i_merge_pe               (merge_valid_i_9_12),
    .data_i_merge_pe                (merge_data_i_9_12),
    .ready_o_merge_pe               (merge_ready_o_9_12),
    .valid_o_merge_pe               (merge_valid_o_9_12),
    .data_o_merge_pe                (merge_data_o_9_12),
    .ready_i_merge_pe               (merge_ready_i_9_12),

    .valid_i_gather_pe              (gather_valid_i_9_12),
    .data_i_gather_pe               (gather_data_i_9_12),
    .ready_o_gather_pe              (gather_ready_o_9_12),
    .valid_o_gather_pe              (gather_valid_o_9_12),
    .data_o_gather_pe               (gather_data_o_9_12),
    .ready_i_gather_pe              (gather_ready_i_9_12),

    .credit_upd                     (credit_upd[9][12])
);


network_interface #(
    .cast_out                       (cast_out_9_13),
    .gather_out                     (gather_out_9_13),
    .cast_sid                       (cast_sid_9_13),
    .gather_sid                     (gather_sid_9_13)
)ni_9_13(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[9][13]),
    .data_i_cast_nw                 (data_o_cast_nw[9][13]),
    .ready_o_cast_nw                (ready_i_cast_nw[9][13]),
    .valid_o_cast_nw                (valid_i_cast_nw[9][13]),
    .data_o_cast_nw                 (data_i_cast_nw[9][13]),
    .ready_i_cast_nw                (ready_o_cast_nw[9][13]),

    .valid_i_gather_nw              (valid_o_gather_nw[9][13]),
    .data_i_gather_nw               (data_o_gather_nw[9][13]),
    .ready_o_gather_nw              (ready_i_gather_nw[9][13]),
    .valid_o_gather_nw              (valid_i_gather_nw[9][13]),
    .data_o_gather_nw               (data_i_gather_nw[9][13]),
    .ready_i_gather_nw              (ready_o_gather_nw[9][13]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[9][13]),
    .data_i_merge_nw                (data_o_merge_nw[9][13]),
    .ready_o_merge_nw               (ready_i_merge_nw[9][13]),
    .valid_o_merge_nw               (valid_i_merge_nw[9][13]),
    .data_o_merge_nw                (data_i_merge_nw[9][13]),
    .ready_i_merge_nw               (ready_o_merge_nw[9][13]),

    .valid_i_cast_pe                (cast_valid_i_9_13),
    .data_i_cast_pe                 (cast_data_i_9_13),
    .ready_o_cast_pe                (cast_ready_o_9_13),
    .valid_o_cast_pe                (cast_valid_o_9_13),
    .data_o_cast_pe                 (cast_data_o_9_13),
    .ready_i_cast_pe                (cast_ready_i_9_13),

    .valid_i_merge_pe               (merge_valid_i_9_13),
    .data_i_merge_pe                (merge_data_i_9_13),
    .ready_o_merge_pe               (merge_ready_o_9_13),
    .valid_o_merge_pe               (merge_valid_o_9_13),
    .data_o_merge_pe                (merge_data_o_9_13),
    .ready_i_merge_pe               (merge_ready_i_9_13),

    .valid_i_gather_pe              (gather_valid_i_9_13),
    .data_i_gather_pe               (gather_data_i_9_13),
    .ready_o_gather_pe              (gather_ready_o_9_13),
    .valid_o_gather_pe              (gather_valid_o_9_13),
    .data_o_gather_pe               (gather_data_o_9_13),
    .ready_i_gather_pe              (gather_ready_i_9_13),

    .credit_upd                     (credit_upd[9][13])
);


network_interface #(
    .cast_out                       (cast_out_9_14),
    .gather_out                     (gather_out_9_14),
    .cast_sid                       (cast_sid_9_14),
    .gather_sid                     (gather_sid_9_14)
)ni_9_14(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[9][14]),
    .data_i_cast_nw                 (data_o_cast_nw[9][14]),
    .ready_o_cast_nw                (ready_i_cast_nw[9][14]),
    .valid_o_cast_nw                (valid_i_cast_nw[9][14]),
    .data_o_cast_nw                 (data_i_cast_nw[9][14]),
    .ready_i_cast_nw                (ready_o_cast_nw[9][14]),

    .valid_i_gather_nw              (valid_o_gather_nw[9][14]),
    .data_i_gather_nw               (data_o_gather_nw[9][14]),
    .ready_o_gather_nw              (ready_i_gather_nw[9][14]),
    .valid_o_gather_nw              (valid_i_gather_nw[9][14]),
    .data_o_gather_nw               (data_i_gather_nw[9][14]),
    .ready_i_gather_nw              (ready_o_gather_nw[9][14]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[9][14]),
    .data_i_merge_nw                (data_o_merge_nw[9][14]),
    .ready_o_merge_nw               (ready_i_merge_nw[9][14]),
    .valid_o_merge_nw               (valid_i_merge_nw[9][14]),
    .data_o_merge_nw                (data_i_merge_nw[9][14]),
    .ready_i_merge_nw               (ready_o_merge_nw[9][14]),

    .valid_i_cast_pe                (cast_valid_i_9_14),
    .data_i_cast_pe                 (cast_data_i_9_14),
    .ready_o_cast_pe                (cast_ready_o_9_14),
    .valid_o_cast_pe                (cast_valid_o_9_14),
    .data_o_cast_pe                 (cast_data_o_9_14),
    .ready_i_cast_pe                (cast_ready_i_9_14),

    .valid_i_merge_pe               (merge_valid_i_9_14),
    .data_i_merge_pe                (merge_data_i_9_14),
    .ready_o_merge_pe               (merge_ready_o_9_14),
    .valid_o_merge_pe               (merge_valid_o_9_14),
    .data_o_merge_pe                (merge_data_o_9_14),
    .ready_i_merge_pe               (merge_ready_i_9_14),

    .valid_i_gather_pe              (gather_valid_i_9_14),
    .data_i_gather_pe               (gather_data_i_9_14),
    .ready_o_gather_pe              (gather_ready_o_9_14),
    .valid_o_gather_pe              (gather_valid_o_9_14),
    .data_o_gather_pe               (gather_data_o_9_14),
    .ready_i_gather_pe              (gather_ready_i_9_14),

    .credit_upd                     (credit_upd[9][14])
);


network_interface #(
    .cast_out                       (cast_out_9_15),
    .gather_out                     (gather_out_9_15),
    .cast_sid                       (cast_sid_9_15),
    .gather_sid                     (gather_sid_9_15)
)ni_9_15(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[9][15]),
    .data_i_cast_nw                 (data_o_cast_nw[9][15]),
    .ready_o_cast_nw                (ready_i_cast_nw[9][15]),
    .valid_o_cast_nw                (valid_i_cast_nw[9][15]),
    .data_o_cast_nw                 (data_i_cast_nw[9][15]),
    .ready_i_cast_nw                (ready_o_cast_nw[9][15]),

    .valid_i_gather_nw              (valid_o_gather_nw[9][15]),
    .data_i_gather_nw               (data_o_gather_nw[9][15]),
    .ready_o_gather_nw              (ready_i_gather_nw[9][15]),
    .valid_o_gather_nw              (valid_i_gather_nw[9][15]),
    .data_o_gather_nw               (data_i_gather_nw[9][15]),
    .ready_i_gather_nw              (ready_o_gather_nw[9][15]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[9][15]),
    .data_i_merge_nw                (data_o_merge_nw[9][15]),
    .ready_o_merge_nw               (ready_i_merge_nw[9][15]),
    .valid_o_merge_nw               (valid_i_merge_nw[9][15]),
    .data_o_merge_nw                (data_i_merge_nw[9][15]),
    .ready_i_merge_nw               (ready_o_merge_nw[9][15]),

    .valid_i_cast_pe                (cast_valid_i_9_15),
    .data_i_cast_pe                 (cast_data_i_9_15),
    .ready_o_cast_pe                (cast_ready_o_9_15),
    .valid_o_cast_pe                (cast_valid_o_9_15),
    .data_o_cast_pe                 (cast_data_o_9_15),
    .ready_i_cast_pe                (cast_ready_i_9_15),

    .valid_i_merge_pe               (merge_valid_i_9_15),
    .data_i_merge_pe                (merge_data_i_9_15),
    .ready_o_merge_pe               (merge_ready_o_9_15),
    .valid_o_merge_pe               (merge_valid_o_9_15),
    .data_o_merge_pe                (merge_data_o_9_15),
    .ready_i_merge_pe               (merge_ready_i_9_15),

    .valid_i_gather_pe              (gather_valid_i_9_15),
    .data_i_gather_pe               (gather_data_i_9_15),
    .ready_o_gather_pe              (gather_ready_o_9_15),
    .valid_o_gather_pe              (gather_valid_o_9_15),
    .data_o_gather_pe               (gather_data_o_9_15),
    .ready_i_gather_pe              (gather_ready_i_9_15),

    .credit_upd                     (credit_upd[9][15])
);


network_interface #(
    .cast_out                       (cast_out_9_16),
    .gather_out                     (gather_out_9_16),
    .cast_sid                       (cast_sid_9_16),
    .gather_sid                     (gather_sid_9_16)
)ni_9_16(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[9][16]),
    .data_i_cast_nw                 (data_o_cast_nw[9][16]),
    .ready_o_cast_nw                (ready_i_cast_nw[9][16]),
    .valid_o_cast_nw                (valid_i_cast_nw[9][16]),
    .data_o_cast_nw                 (data_i_cast_nw[9][16]),
    .ready_i_cast_nw                (ready_o_cast_nw[9][16]),

    .valid_i_gather_nw              (valid_o_gather_nw[9][16]),
    .data_i_gather_nw               (data_o_gather_nw[9][16]),
    .ready_o_gather_nw              (ready_i_gather_nw[9][16]),
    .valid_o_gather_nw              (valid_i_gather_nw[9][16]),
    .data_o_gather_nw               (data_i_gather_nw[9][16]),
    .ready_i_gather_nw              (ready_o_gather_nw[9][16]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[9][16]),
    .data_i_merge_nw                (data_o_merge_nw[9][16]),
    .ready_o_merge_nw               (ready_i_merge_nw[9][16]),
    .valid_o_merge_nw               (valid_i_merge_nw[9][16]),
    .data_o_merge_nw                (data_i_merge_nw[9][16]),
    .ready_i_merge_nw               (ready_o_merge_nw[9][16]),

    .valid_i_cast_pe                (cast_valid_i_9_16),
    .data_i_cast_pe                 (cast_data_i_9_16),
    .ready_o_cast_pe                (cast_ready_o_9_16),
    .valid_o_cast_pe                (cast_valid_o_9_16),
    .data_o_cast_pe                 (cast_data_o_9_16),
    .ready_i_cast_pe                (cast_ready_i_9_16),

    .valid_i_merge_pe               (merge_valid_i_9_16),
    .data_i_merge_pe                (merge_data_i_9_16),
    .ready_o_merge_pe               (merge_ready_o_9_16),
    .valid_o_merge_pe               (merge_valid_o_9_16),
    .data_o_merge_pe                (merge_data_o_9_16),
    .ready_i_merge_pe               (merge_ready_i_9_16),

    .valid_i_gather_pe              (gather_valid_i_9_16),
    .data_i_gather_pe               (gather_data_i_9_16),
    .ready_o_gather_pe              (gather_ready_o_9_16),
    .valid_o_gather_pe              (gather_valid_o_9_16),
    .data_o_gather_pe               (gather_data_o_9_16),
    .ready_i_gather_pe              (gather_ready_i_9_16),

    .credit_upd                     (credit_upd[9][16])
);


network_interface #(
    .cast_out                       (cast_out_9_17),
    .gather_out                     (gather_out_9_17),
    .cast_sid                       (cast_sid_9_17),
    .gather_sid                     (gather_sid_9_17)
)ni_9_17(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[9][17]),
    .data_i_cast_nw                 (data_o_cast_nw[9][17]),
    .ready_o_cast_nw                (ready_i_cast_nw[9][17]),
    .valid_o_cast_nw                (valid_i_cast_nw[9][17]),
    .data_o_cast_nw                 (data_i_cast_nw[9][17]),
    .ready_i_cast_nw                (ready_o_cast_nw[9][17]),

    .valid_i_gather_nw              (valid_o_gather_nw[9][17]),
    .data_i_gather_nw               (data_o_gather_nw[9][17]),
    .ready_o_gather_nw              (ready_i_gather_nw[9][17]),
    .valid_o_gather_nw              (valid_i_gather_nw[9][17]),
    .data_o_gather_nw               (data_i_gather_nw[9][17]),
    .ready_i_gather_nw              (ready_o_gather_nw[9][17]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[9][17]),
    .data_i_merge_nw                (data_o_merge_nw[9][17]),
    .ready_o_merge_nw               (ready_i_merge_nw[9][17]),
    .valid_o_merge_nw               (valid_i_merge_nw[9][17]),
    .data_o_merge_nw                (data_i_merge_nw[9][17]),
    .ready_i_merge_nw               (ready_o_merge_nw[9][17]),

    .valid_i_cast_pe                (cast_valid_i_9_17),
    .data_i_cast_pe                 (cast_data_i_9_17),
    .ready_o_cast_pe                (cast_ready_o_9_17),
    .valid_o_cast_pe                (cast_valid_o_9_17),
    .data_o_cast_pe                 (cast_data_o_9_17),
    .ready_i_cast_pe                (cast_ready_i_9_17),

    .valid_i_merge_pe               (merge_valid_i_9_17),
    .data_i_merge_pe                (merge_data_i_9_17),
    .ready_o_merge_pe               (merge_ready_o_9_17),
    .valid_o_merge_pe               (merge_valid_o_9_17),
    .data_o_merge_pe                (merge_data_o_9_17),
    .ready_i_merge_pe               (merge_ready_i_9_17),

    .valid_i_gather_pe              (gather_valid_i_9_17),
    .data_i_gather_pe               (gather_data_i_9_17),
    .ready_o_gather_pe              (gather_ready_o_9_17),
    .valid_o_gather_pe              (gather_valid_o_9_17),
    .data_o_gather_pe               (gather_data_o_9_17),
    .ready_i_gather_pe              (gather_ready_i_9_17),

    .credit_upd                     (credit_upd[9][17])
);


network_interface #(
    .cast_out                       (cast_out_9_18),
    .gather_out                     (gather_out_9_18),
    .cast_sid                       (cast_sid_9_18),
    .gather_sid                     (gather_sid_9_18)
)ni_9_18(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[9][18]),
    .data_i_cast_nw                 (data_o_cast_nw[9][18]),
    .ready_o_cast_nw                (ready_i_cast_nw[9][18]),
    .valid_o_cast_nw                (valid_i_cast_nw[9][18]),
    .data_o_cast_nw                 (data_i_cast_nw[9][18]),
    .ready_i_cast_nw                (ready_o_cast_nw[9][18]),

    .valid_i_gather_nw              (valid_o_gather_nw[9][18]),
    .data_i_gather_nw               (data_o_gather_nw[9][18]),
    .ready_o_gather_nw              (ready_i_gather_nw[9][18]),
    .valid_o_gather_nw              (valid_i_gather_nw[9][18]),
    .data_o_gather_nw               (data_i_gather_nw[9][18]),
    .ready_i_gather_nw              (ready_o_gather_nw[9][18]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[9][18]),
    .data_i_merge_nw                (data_o_merge_nw[9][18]),
    .ready_o_merge_nw               (ready_i_merge_nw[9][18]),
    .valid_o_merge_nw               (valid_i_merge_nw[9][18]),
    .data_o_merge_nw                (data_i_merge_nw[9][18]),
    .ready_i_merge_nw               (ready_o_merge_nw[9][18]),

    .valid_i_cast_pe                (cast_valid_i_9_18),
    .data_i_cast_pe                 (cast_data_i_9_18),
    .ready_o_cast_pe                (cast_ready_o_9_18),
    .valid_o_cast_pe                (cast_valid_o_9_18),
    .data_o_cast_pe                 (cast_data_o_9_18),
    .ready_i_cast_pe                (cast_ready_i_9_18),

    .valid_i_merge_pe               (merge_valid_i_9_18),
    .data_i_merge_pe                (merge_data_i_9_18),
    .ready_o_merge_pe               (merge_ready_o_9_18),
    .valid_o_merge_pe               (merge_valid_o_9_18),
    .data_o_merge_pe                (merge_data_o_9_18),
    .ready_i_merge_pe               (merge_ready_i_9_18),

    .valid_i_gather_pe              (gather_valid_i_9_18),
    .data_i_gather_pe               (gather_data_i_9_18),
    .ready_o_gather_pe              (gather_ready_o_9_18),
    .valid_o_gather_pe              (gather_valid_o_9_18),
    .data_o_gather_pe               (gather_data_o_9_18),
    .ready_i_gather_pe              (gather_ready_i_9_18),

    .credit_upd                     (credit_upd[9][18])
);


network_interface #(
    .cast_out                       (cast_out_9_19),
    .gather_out                     (gather_out_9_19),
    .cast_sid                       (cast_sid_9_19),
    .gather_sid                     (gather_sid_9_19)
)ni_9_19(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[9][19]),
    .data_i_cast_nw                 (data_o_cast_nw[9][19]),
    .ready_o_cast_nw                (ready_i_cast_nw[9][19]),
    .valid_o_cast_nw                (valid_i_cast_nw[9][19]),
    .data_o_cast_nw                 (data_i_cast_nw[9][19]),
    .ready_i_cast_nw                (ready_o_cast_nw[9][19]),

    .valid_i_gather_nw              (valid_o_gather_nw[9][19]),
    .data_i_gather_nw               (data_o_gather_nw[9][19]),
    .ready_o_gather_nw              (ready_i_gather_nw[9][19]),
    .valid_o_gather_nw              (valid_i_gather_nw[9][19]),
    .data_o_gather_nw               (data_i_gather_nw[9][19]),
    .ready_i_gather_nw              (ready_o_gather_nw[9][19]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[9][19]),
    .data_i_merge_nw                (data_o_merge_nw[9][19]),
    .ready_o_merge_nw               (ready_i_merge_nw[9][19]),
    .valid_o_merge_nw               (valid_i_merge_nw[9][19]),
    .data_o_merge_nw                (data_i_merge_nw[9][19]),
    .ready_i_merge_nw               (ready_o_merge_nw[9][19]),

    .valid_i_cast_pe                (cast_valid_i_9_19),
    .data_i_cast_pe                 (cast_data_i_9_19),
    .ready_o_cast_pe                (cast_ready_o_9_19),
    .valid_o_cast_pe                (cast_valid_o_9_19),
    .data_o_cast_pe                 (cast_data_o_9_19),
    .ready_i_cast_pe                (cast_ready_i_9_19),

    .valid_i_merge_pe               (merge_valid_i_9_19),
    .data_i_merge_pe                (merge_data_i_9_19),
    .ready_o_merge_pe               (merge_ready_o_9_19),
    .valid_o_merge_pe               (merge_valid_o_9_19),
    .data_o_merge_pe                (merge_data_o_9_19),
    .ready_i_merge_pe               (merge_ready_i_9_19),

    .valid_i_gather_pe              (gather_valid_i_9_19),
    .data_i_gather_pe               (gather_data_i_9_19),
    .ready_o_gather_pe              (gather_ready_o_9_19),
    .valid_o_gather_pe              (gather_valid_o_9_19),
    .data_o_gather_pe               (gather_data_o_9_19),
    .ready_i_gather_pe              (gather_ready_i_9_19),

    .credit_upd                     (credit_upd[9][19])
);


network_interface #(
    .cast_out                       (cast_out_9_20),
    .gather_out                     (gather_out_9_20),
    .cast_sid                       (cast_sid_9_20),
    .gather_sid                     (gather_sid_9_20)
)ni_9_20(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[9][20]),
    .data_i_cast_nw                 (data_o_cast_nw[9][20]),
    .ready_o_cast_nw                (ready_i_cast_nw[9][20]),
    .valid_o_cast_nw                (valid_i_cast_nw[9][20]),
    .data_o_cast_nw                 (data_i_cast_nw[9][20]),
    .ready_i_cast_nw                (ready_o_cast_nw[9][20]),

    .valid_i_gather_nw              (valid_o_gather_nw[9][20]),
    .data_i_gather_nw               (data_o_gather_nw[9][20]),
    .ready_o_gather_nw              (ready_i_gather_nw[9][20]),
    .valid_o_gather_nw              (valid_i_gather_nw[9][20]),
    .data_o_gather_nw               (data_i_gather_nw[9][20]),
    .ready_i_gather_nw              (ready_o_gather_nw[9][20]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[9][20]),
    .data_i_merge_nw                (data_o_merge_nw[9][20]),
    .ready_o_merge_nw               (ready_i_merge_nw[9][20]),
    .valid_o_merge_nw               (valid_i_merge_nw[9][20]),
    .data_o_merge_nw                (data_i_merge_nw[9][20]),
    .ready_i_merge_nw               (ready_o_merge_nw[9][20]),

    .valid_i_cast_pe                (cast_valid_i_9_20),
    .data_i_cast_pe                 (cast_data_i_9_20),
    .ready_o_cast_pe                (cast_ready_o_9_20),
    .valid_o_cast_pe                (cast_valid_o_9_20),
    .data_o_cast_pe                 (cast_data_o_9_20),
    .ready_i_cast_pe                (cast_ready_i_9_20),

    .valid_i_merge_pe               (merge_valid_i_9_20),
    .data_i_merge_pe                (merge_data_i_9_20),
    .ready_o_merge_pe               (merge_ready_o_9_20),
    .valid_o_merge_pe               (merge_valid_o_9_20),
    .data_o_merge_pe                (merge_data_o_9_20),
    .ready_i_merge_pe               (merge_ready_i_9_20),

    .valid_i_gather_pe              (gather_valid_i_9_20),
    .data_i_gather_pe               (gather_data_i_9_20),
    .ready_o_gather_pe              (gather_ready_o_9_20),
    .valid_o_gather_pe              (gather_valid_o_9_20),
    .data_o_gather_pe               (gather_data_o_9_20),
    .ready_i_gather_pe              (gather_ready_i_9_20),

    .credit_upd                     (credit_upd[9][20])
);


network_interface #(
    .cast_out                       (cast_out_9_21),
    .gather_out                     (gather_out_9_21),
    .cast_sid                       (cast_sid_9_21),
    .gather_sid                     (gather_sid_9_21)
)ni_9_21(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[9][21]),
    .data_i_cast_nw                 (data_o_cast_nw[9][21]),
    .ready_o_cast_nw                (ready_i_cast_nw[9][21]),
    .valid_o_cast_nw                (valid_i_cast_nw[9][21]),
    .data_o_cast_nw                 (data_i_cast_nw[9][21]),
    .ready_i_cast_nw                (ready_o_cast_nw[9][21]),

    .valid_i_gather_nw              (valid_o_gather_nw[9][21]),
    .data_i_gather_nw               (data_o_gather_nw[9][21]),
    .ready_o_gather_nw              (ready_i_gather_nw[9][21]),
    .valid_o_gather_nw              (valid_i_gather_nw[9][21]),
    .data_o_gather_nw               (data_i_gather_nw[9][21]),
    .ready_i_gather_nw              (ready_o_gather_nw[9][21]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[9][21]),
    .data_i_merge_nw                (data_o_merge_nw[9][21]),
    .ready_o_merge_nw               (ready_i_merge_nw[9][21]),
    .valid_o_merge_nw               (valid_i_merge_nw[9][21]),
    .data_o_merge_nw                (data_i_merge_nw[9][21]),
    .ready_i_merge_nw               (ready_o_merge_nw[9][21]),

    .valid_i_cast_pe                (cast_valid_i_9_21),
    .data_i_cast_pe                 (cast_data_i_9_21),
    .ready_o_cast_pe                (cast_ready_o_9_21),
    .valid_o_cast_pe                (cast_valid_o_9_21),
    .data_o_cast_pe                 (cast_data_o_9_21),
    .ready_i_cast_pe                (cast_ready_i_9_21),

    .valid_i_merge_pe               (merge_valid_i_9_21),
    .data_i_merge_pe                (merge_data_i_9_21),
    .ready_o_merge_pe               (merge_ready_o_9_21),
    .valid_o_merge_pe               (merge_valid_o_9_21),
    .data_o_merge_pe                (merge_data_o_9_21),
    .ready_i_merge_pe               (merge_ready_i_9_21),

    .valid_i_gather_pe              (gather_valid_i_9_21),
    .data_i_gather_pe               (gather_data_i_9_21),
    .ready_o_gather_pe              (gather_ready_o_9_21),
    .valid_o_gather_pe              (gather_valid_o_9_21),
    .data_o_gather_pe               (gather_data_o_9_21),
    .ready_i_gather_pe              (gather_ready_i_9_21),

    .credit_upd                     (credit_upd[9][21])
);


network_interface #(
    .cast_out                       (cast_out_9_22),
    .gather_out                     (gather_out_9_22),
    .cast_sid                       (cast_sid_9_22),
    .gather_sid                     (gather_sid_9_22)
)ni_9_22(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[9][22]),
    .data_i_cast_nw                 (data_o_cast_nw[9][22]),
    .ready_o_cast_nw                (ready_i_cast_nw[9][22]),
    .valid_o_cast_nw                (valid_i_cast_nw[9][22]),
    .data_o_cast_nw                 (data_i_cast_nw[9][22]),
    .ready_i_cast_nw                (ready_o_cast_nw[9][22]),

    .valid_i_gather_nw              (valid_o_gather_nw[9][22]),
    .data_i_gather_nw               (data_o_gather_nw[9][22]),
    .ready_o_gather_nw              (ready_i_gather_nw[9][22]),
    .valid_o_gather_nw              (valid_i_gather_nw[9][22]),
    .data_o_gather_nw               (data_i_gather_nw[9][22]),
    .ready_i_gather_nw              (ready_o_gather_nw[9][22]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[9][22]),
    .data_i_merge_nw                (data_o_merge_nw[9][22]),
    .ready_o_merge_nw               (ready_i_merge_nw[9][22]),
    .valid_o_merge_nw               (valid_i_merge_nw[9][22]),
    .data_o_merge_nw                (data_i_merge_nw[9][22]),
    .ready_i_merge_nw               (ready_o_merge_nw[9][22]),

    .valid_i_cast_pe                (cast_valid_i_9_22),
    .data_i_cast_pe                 (cast_data_i_9_22),
    .ready_o_cast_pe                (cast_ready_o_9_22),
    .valid_o_cast_pe                (cast_valid_o_9_22),
    .data_o_cast_pe                 (cast_data_o_9_22),
    .ready_i_cast_pe                (cast_ready_i_9_22),

    .valid_i_merge_pe               (merge_valid_i_9_22),
    .data_i_merge_pe                (merge_data_i_9_22),
    .ready_o_merge_pe               (merge_ready_o_9_22),
    .valid_o_merge_pe               (merge_valid_o_9_22),
    .data_o_merge_pe                (merge_data_o_9_22),
    .ready_i_merge_pe               (merge_ready_i_9_22),

    .valid_i_gather_pe              (gather_valid_i_9_22),
    .data_i_gather_pe               (gather_data_i_9_22),
    .ready_o_gather_pe              (gather_ready_o_9_22),
    .valid_o_gather_pe              (gather_valid_o_9_22),
    .data_o_gather_pe               (gather_data_o_9_22),
    .ready_i_gather_pe              (gather_ready_i_9_22),

    .credit_upd                     (credit_upd[9][22])
);


network_interface #(
    .cast_out                       (cast_out_9_23),
    .gather_out                     (gather_out_9_23),
    .cast_sid                       (cast_sid_9_23),
    .gather_sid                     (gather_sid_9_23)
)ni_9_23(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[9][23]),
    .data_i_cast_nw                 (data_o_cast_nw[9][23]),
    .ready_o_cast_nw                (ready_i_cast_nw[9][23]),
    .valid_o_cast_nw                (valid_i_cast_nw[9][23]),
    .data_o_cast_nw                 (data_i_cast_nw[9][23]),
    .ready_i_cast_nw                (ready_o_cast_nw[9][23]),

    .valid_i_gather_nw              (valid_o_gather_nw[9][23]),
    .data_i_gather_nw               (data_o_gather_nw[9][23]),
    .ready_o_gather_nw              (ready_i_gather_nw[9][23]),
    .valid_o_gather_nw              (valid_i_gather_nw[9][23]),
    .data_o_gather_nw               (data_i_gather_nw[9][23]),
    .ready_i_gather_nw              (ready_o_gather_nw[9][23]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[9][23]),
    .data_i_merge_nw                (data_o_merge_nw[9][23]),
    .ready_o_merge_nw               (ready_i_merge_nw[9][23]),
    .valid_o_merge_nw               (valid_i_merge_nw[9][23]),
    .data_o_merge_nw                (data_i_merge_nw[9][23]),
    .ready_i_merge_nw               (ready_o_merge_nw[9][23]),

    .valid_i_cast_pe                (cast_valid_i_9_23),
    .data_i_cast_pe                 (cast_data_i_9_23),
    .ready_o_cast_pe                (cast_ready_o_9_23),
    .valid_o_cast_pe                (cast_valid_o_9_23),
    .data_o_cast_pe                 (cast_data_o_9_23),
    .ready_i_cast_pe                (cast_ready_i_9_23),

    .valid_i_merge_pe               (merge_valid_i_9_23),
    .data_i_merge_pe                (merge_data_i_9_23),
    .ready_o_merge_pe               (merge_ready_o_9_23),
    .valid_o_merge_pe               (merge_valid_o_9_23),
    .data_o_merge_pe                (merge_data_o_9_23),
    .ready_i_merge_pe               (merge_ready_i_9_23),

    .valid_i_gather_pe              (gather_valid_i_9_23),
    .data_i_gather_pe               (gather_data_i_9_23),
    .ready_o_gather_pe              (gather_ready_o_9_23),
    .valid_o_gather_pe              (gather_valid_o_9_23),
    .data_o_gather_pe               (gather_data_o_9_23),
    .ready_i_gather_pe              (gather_ready_i_9_23),

    .credit_upd                     (credit_upd[9][23])
);


network_interface #(
    .cast_out                       (cast_out_9_24),
    .gather_out                     (gather_out_9_24),
    .cast_sid                       (cast_sid_9_24),
    .gather_sid                     (gather_sid_9_24)
)ni_9_24(
    .clk                            (clk),
    .rstn                           (rstn),

    .valid_i_cast_nw                (valid_o_cast_nw[9][24]),
    .data_i_cast_nw                 (data_o_cast_nw[9][24]),
    .ready_o_cast_nw                (ready_i_cast_nw[9][24]),
    .valid_o_cast_nw                (valid_i_cast_nw[9][24]),
    .data_o_cast_nw                 (data_i_cast_nw[9][24]),
    .ready_i_cast_nw                (ready_o_cast_nw[9][24]),

    .valid_i_gather_nw              (valid_o_gather_nw[9][24]),
    .data_i_gather_nw               (data_o_gather_nw[9][24]),
    .ready_o_gather_nw              (ready_i_gather_nw[9][24]),
    .valid_o_gather_nw              (valid_i_gather_nw[9][24]),
    .data_o_gather_nw               (data_i_gather_nw[9][24]),
    .ready_i_gather_nw              (ready_o_gather_nw[9][24]),
    
    .valid_i_merge_nw               (valid_o_merge_nw[9][24]),
    .data_i_merge_nw                (data_o_merge_nw[9][24]),
    .ready_o_merge_nw               (ready_i_merge_nw[9][24]),
    .valid_o_merge_nw               (valid_i_merge_nw[9][24]),
    .data_o_merge_nw                (data_i_merge_nw[9][24]),
    .ready_i_merge_nw               (ready_o_merge_nw[9][24]),

    .valid_i_cast_pe                (cast_valid_i_9_24),
    .data_i_cast_pe                 (cast_data_i_9_24),
    .ready_o_cast_pe                (cast_ready_o_9_24),
    .valid_o_cast_pe                (cast_valid_o_9_24),
    .data_o_cast_pe                 (cast_data_o_9_24),
    .ready_i_cast_pe                (cast_ready_i_9_24),

    .valid_i_merge_pe               (merge_valid_i_9_24),
    .data_i_merge_pe                (merge_data_i_9_24),
    .ready_o_merge_pe               (merge_ready_o_9_24),
    .valid_o_merge_pe               (merge_valid_o_9_24),
    .data_o_merge_pe                (merge_data_o_9_24),
    .ready_i_merge_pe               (merge_ready_i_9_24),

    .valid_i_gather_pe              (gather_valid_i_9_24),
    .data_i_gather_pe               (gather_data_i_9_24),
    .ready_o_gather_pe              (gather_ready_o_9_24),
    .valid_o_gather_pe              (gather_valid_o_9_24),
    .data_o_gather_pe               (gather_data_o_9_24),
    .ready_i_gather_pe              (gather_ready_i_9_24),

    .credit_upd                     (credit_upd[9][24])
);

endmodule
