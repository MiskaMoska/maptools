
`ifndef __NETWORK_CONFIG_SVH_
`define __NETWORK_CONFIG_SVH_
    
localparam cast_out_0_0 = 1;
localparam merge_out_0_0 = 0;
localparam gather_out_0_0 = 0;
localparam merge_in_0_0 = 0;
localparam gather_in_0_0 = 0;
localparam cast_sid_0_0 = 1;
localparam gather_sid_0_0 = 0;

localparam cast_out_0_1 = 1;
localparam merge_out_0_1 = 0;
localparam gather_out_0_1 = 0;
localparam merge_in_0_1 = 0;
localparam gather_in_0_1 = 0;
localparam cast_sid_0_1 = 16;
localparam gather_sid_0_1 = 0;

localparam cast_out_0_2 = 1;
localparam merge_out_0_2 = 0;
localparam gather_out_0_2 = 1;
localparam merge_in_0_2 = 0;
localparam gather_in_0_2 = 1;
localparam cast_sid_0_2 = 17;
localparam gather_sid_0_2 = 8;

localparam cast_out_0_3 = 0;
localparam merge_out_0_3 = 0;
localparam gather_out_0_3 = 1;
localparam merge_in_0_3 = 1;
localparam gather_in_0_3 = 0;
localparam cast_sid_0_3 = 0;
localparam gather_sid_0_3 = 18;

localparam cast_out_0_4 = 0;
localparam merge_out_0_4 = 1;
localparam gather_out_0_4 = 0;
localparam merge_in_0_4 = 0;
localparam gather_in_0_4 = 0;
localparam cast_sid_0_4 = 0;
localparam gather_sid_0_4 = 0;

localparam cast_out_0_5 = 0;
localparam merge_out_0_5 = 1;
localparam gather_out_0_5 = 0;
localparam merge_in_0_5 = 0;
localparam gather_in_0_5 = 0;
localparam cast_sid_0_5 = 0;
localparam gather_sid_0_5 = 0;

localparam cast_out_0_6 = 0;
localparam merge_out_0_6 = 1;
localparam gather_out_0_6 = 0;
localparam merge_in_0_6 = 0;
localparam gather_in_0_6 = 0;
localparam cast_sid_0_6 = 0;
localparam gather_sid_0_6 = 0;

localparam cast_out_0_7 = 0;
localparam merge_out_0_7 = 1;
localparam gather_out_0_7 = 0;
localparam merge_in_0_7 = 0;
localparam gather_in_0_7 = 0;
localparam cast_sid_0_7 = 0;
localparam gather_sid_0_7 = 0;

localparam cast_out_0_8 = 0;
localparam merge_out_0_8 = 1;
localparam gather_out_0_8 = 0;
localparam merge_in_0_8 = 0;
localparam gather_in_0_8 = 0;
localparam cast_sid_0_8 = 0;
localparam gather_sid_0_8 = 0;

localparam cast_out_0_9 = 0;
localparam merge_out_0_9 = 1;
localparam gather_out_0_9 = 0;
localparam merge_in_0_9 = 0;
localparam gather_in_0_9 = 0;
localparam cast_sid_0_9 = 0;
localparam gather_sid_0_9 = 0;

localparam cast_out_0_10 = 0;
localparam merge_out_0_10 = 1;
localparam gather_out_0_10 = 0;
localparam merge_in_0_10 = 0;
localparam gather_in_0_10 = 0;
localparam cast_sid_0_10 = 0;
localparam gather_sid_0_10 = 0;

localparam cast_out_0_11 = 0;
localparam merge_out_0_11 = 1;
localparam gather_out_0_11 = 0;
localparam merge_in_0_11 = 0;
localparam gather_in_0_11 = 0;
localparam cast_sid_0_11 = 0;
localparam gather_sid_0_11 = 0;

localparam cast_out_0_12 = 0;
localparam merge_out_0_12 = 1;
localparam gather_out_0_12 = 0;
localparam merge_in_0_12 = 0;
localparam gather_in_0_12 = 0;
localparam cast_sid_0_12 = 0;
localparam gather_sid_0_12 = 0;

localparam cast_out_0_13 = 0;
localparam merge_out_0_13 = 1;
localparam gather_out_0_13 = 0;
localparam merge_in_0_13 = 0;
localparam gather_in_0_13 = 0;
localparam cast_sid_0_13 = 0;
localparam gather_sid_0_13 = 0;

localparam cast_out_0_14 = 0;
localparam merge_out_0_14 = 1;
localparam gather_out_0_14 = 0;
localparam merge_in_0_14 = 0;
localparam gather_in_0_14 = 0;
localparam cast_sid_0_14 = 0;
localparam gather_sid_0_14 = 0;

localparam cast_out_0_15 = 0;
localparam merge_out_0_15 = 1;
localparam gather_out_0_15 = 0;
localparam merge_in_0_15 = 0;
localparam gather_in_0_15 = 0;
localparam cast_sid_0_15 = 0;
localparam gather_sid_0_15 = 0;

localparam cast_out_0_16 = 0;
localparam merge_out_0_16 = 1;
localparam gather_out_0_16 = 0;
localparam merge_in_0_16 = 0;
localparam gather_in_0_16 = 0;
localparam cast_sid_0_16 = 0;
localparam gather_sid_0_16 = 0;

localparam cast_out_0_17 = 0;
localparam merge_out_0_17 = 1;
localparam gather_out_0_17 = 0;
localparam merge_in_0_17 = 0;
localparam gather_in_0_17 = 0;
localparam cast_sid_0_17 = 0;
localparam gather_sid_0_17 = 0;

localparam cast_out_0_18 = 0;
localparam merge_out_0_18 = 1;
localparam gather_out_0_18 = 0;
localparam merge_in_0_18 = 0;
localparam gather_in_0_18 = 0;
localparam cast_sid_0_18 = 0;
localparam gather_sid_0_18 = 0;

localparam cast_out_0_19 = 0;
localparam merge_out_0_19 = 1;
localparam gather_out_0_19 = 0;
localparam merge_in_0_19 = 0;
localparam gather_in_0_19 = 0;
localparam cast_sid_0_19 = 0;
localparam gather_sid_0_19 = 0;

localparam cast_out_0_20 = 0;
localparam merge_out_0_20 = 1;
localparam gather_out_0_20 = 0;
localparam merge_in_0_20 = 0;
localparam gather_in_0_20 = 0;
localparam cast_sid_0_20 = 0;
localparam gather_sid_0_20 = 0;

localparam cast_out_0_21 = 0;
localparam merge_out_0_21 = 1;
localparam gather_out_0_21 = 0;
localparam merge_in_0_21 = 0;
localparam gather_in_0_21 = 0;
localparam cast_sid_0_21 = 0;
localparam gather_sid_0_21 = 0;

localparam cast_out_0_22 = 0;
localparam merge_out_0_22 = 1;
localparam gather_out_0_22 = 0;
localparam merge_in_0_22 = 0;
localparam gather_in_0_22 = 0;
localparam cast_sid_0_22 = 0;
localparam gather_sid_0_22 = 0;

localparam cast_out_0_23 = 1;
localparam merge_out_0_23 = 0;
localparam gather_out_0_23 = 0;
localparam merge_in_0_23 = 1;
localparam gather_in_0_23 = 1;
localparam cast_sid_0_23 = 1022;
localparam gather_sid_0_23 = 0;

localparam cast_out_0_24 = 0;
localparam merge_out_0_24 = 1;
localparam gather_out_0_24 = 0;
localparam merge_in_0_24 = 0;
localparam gather_in_0_24 = 0;
localparam cast_sid_0_24 = 0;
localparam gather_sid_0_24 = 0;

localparam cast_out_1_0 = 1;
localparam merge_out_1_0 = 0;
localparam gather_out_1_0 = 0;
localparam merge_in_1_0 = 0;
localparam gather_in_1_0 = 0;
localparam cast_sid_1_0 = 2;
localparam gather_sid_1_0 = 0;

localparam cast_out_1_1 = 0;
localparam merge_out_1_1 = 1;
localparam gather_out_1_1 = 0;
localparam merge_in_1_1 = 0;
localparam gather_in_1_1 = 0;
localparam cast_sid_1_1 = 0;
localparam gather_sid_1_1 = 0;

localparam cast_out_1_2 = 1;
localparam merge_out_1_2 = 0;
localparam gather_out_1_2 = 1;
localparam merge_in_1_2 = 0;
localparam gather_in_1_2 = 1;
localparam cast_sid_1_2 = 18;
localparam gather_sid_1_2 = 9;

localparam cast_out_1_3 = 0;
localparam merge_out_1_3 = 1;
localparam gather_out_1_3 = 0;
localparam merge_in_1_3 = 0;
localparam gather_in_1_3 = 0;
localparam cast_sid_1_3 = 0;
localparam gather_sid_1_3 = 0;

localparam cast_out_1_4 = 0;
localparam merge_out_1_4 = 0;
localparam gather_out_1_4 = 1;
localparam merge_in_1_4 = 1;
localparam gather_in_1_4 = 0;
localparam cast_sid_1_4 = 0;
localparam gather_sid_1_4 = 19;

localparam cast_out_1_5 = 0;
localparam merge_out_1_5 = 1;
localparam gather_out_1_5 = 0;
localparam merge_in_1_5 = 0;
localparam gather_in_1_5 = 0;
localparam cast_sid_1_5 = 0;
localparam gather_sid_1_5 = 0;

localparam cast_out_1_6 = 1;
localparam merge_out_1_6 = 0;
localparam gather_out_1_6 = 0;
localparam merge_in_1_6 = 1;
localparam gather_in_1_6 = 0;
localparam cast_sid_1_6 = 39;
localparam gather_sid_1_6 = 0;

localparam cast_out_1_7 = 0;
localparam merge_out_1_7 = 1;
localparam gather_out_1_7 = 0;
localparam merge_in_1_7 = 0;
localparam gather_in_1_7 = 0;
localparam cast_sid_1_7 = 0;
localparam gather_sid_1_7 = 0;

localparam cast_out_1_8 = 1;
localparam merge_out_1_8 = 0;
localparam gather_out_1_8 = 0;
localparam merge_in_1_8 = 1;
localparam gather_in_1_8 = 0;
localparam cast_sid_1_8 = 51;
localparam gather_sid_1_8 = 0;

localparam cast_out_1_9 = 0;
localparam merge_out_1_9 = 1;
localparam gather_out_1_9 = 0;
localparam merge_in_1_9 = 0;
localparam gather_in_1_9 = 0;
localparam cast_sid_1_9 = 0;
localparam gather_sid_1_9 = 0;

localparam cast_out_1_10 = 1;
localparam merge_out_1_10 = 0;
localparam gather_out_1_10 = 0;
localparam merge_in_1_10 = 1;
localparam gather_in_1_10 = 0;
localparam cast_sid_1_10 = 63;
localparam gather_sid_1_10 = 0;

localparam cast_out_1_11 = 0;
localparam merge_out_1_11 = 1;
localparam gather_out_1_11 = 0;
localparam merge_in_1_11 = 0;
localparam gather_in_1_11 = 0;
localparam cast_sid_1_11 = 0;
localparam gather_sid_1_11 = 0;

localparam cast_out_1_12 = 0;
localparam merge_out_1_12 = 0;
localparam gather_out_1_12 = 1;
localparam merge_in_1_12 = 1;
localparam gather_in_1_12 = 0;
localparam cast_sid_1_12 = 0;
localparam gather_sid_1_12 = 47;

localparam cast_out_1_13 = 0;
localparam merge_out_1_13 = 1;
localparam gather_out_1_13 = 0;
localparam merge_in_1_13 = 0;
localparam gather_in_1_13 = 0;
localparam cast_sid_1_13 = 0;
localparam gather_sid_1_13 = 0;

localparam cast_out_1_14 = 1;
localparam merge_out_1_14 = 0;
localparam gather_out_1_14 = 0;
localparam merge_in_1_14 = 1;
localparam gather_in_1_14 = 0;
localparam cast_sid_1_14 = 65;
localparam gather_sid_1_14 = 0;

localparam cast_out_1_15 = 1;
localparam merge_out_1_15 = 0;
localparam gather_out_1_15 = 1;
localparam merge_in_1_15 = 1;
localparam gather_in_1_15 = 1;
localparam cast_sid_1_15 = 73;
localparam gather_sid_1_15 = 42;

localparam cast_out_1_16 = 1;
localparam merge_out_1_16 = 0;
localparam gather_out_1_16 = 1;
localparam merge_in_1_16 = 1;
localparam gather_in_1_16 = 1;
localparam cast_sid_1_16 = 74;
localparam gather_sid_1_16 = 43;

localparam cast_out_1_17 = 0;
localparam merge_out_1_17 = 1;
localparam gather_out_1_17 = 0;
localparam merge_in_1_17 = 0;
localparam gather_in_1_17 = 0;
localparam cast_sid_1_17 = 0;
localparam gather_sid_1_17 = 0;

localparam cast_out_1_18 = 1;
localparam merge_out_1_18 = 0;
localparam gather_out_1_18 = 0;
localparam merge_in_1_18 = 1;
localparam gather_in_1_18 = 0;
localparam cast_sid_1_18 = 77;
localparam gather_sid_1_18 = 0;

localparam cast_out_1_19 = 1;
localparam merge_out_1_19 = 0;
localparam gather_out_1_19 = 1;
localparam merge_in_1_19 = 1;
localparam gather_in_1_19 = 1;
localparam cast_sid_1_19 = 85;
localparam gather_sid_1_19 = 58;

localparam cast_out_1_20 = 1;
localparam merge_out_1_20 = 0;
localparam gather_out_1_20 = 1;
localparam merge_in_1_20 = 1;
localparam gather_in_1_20 = 1;
localparam cast_sid_1_20 = 86;
localparam gather_sid_1_20 = 59;

localparam cast_out_1_21 = 0;
localparam merge_out_1_21 = 1;
localparam gather_out_1_21 = 0;
localparam merge_in_1_21 = 0;
localparam gather_in_1_21 = 0;
localparam cast_sid_1_21 = 0;
localparam gather_sid_1_21 = 0;

localparam cast_out_1_22 = 1;
localparam merge_out_1_22 = 0;
localparam gather_out_1_22 = 0;
localparam merge_in_1_22 = 1;
localparam gather_in_1_22 = 0;
localparam cast_sid_1_22 = 89;
localparam gather_sid_1_22 = 0;

localparam cast_out_1_23 = 0;
localparam merge_out_1_23 = 1;
localparam gather_out_1_23 = 0;
localparam merge_in_1_23 = 0;
localparam gather_in_1_23 = 0;
localparam cast_sid_1_23 = 0;
localparam gather_sid_1_23 = 0;

localparam cast_out_1_24 = 1;
localparam merge_out_1_24 = 0;
localparam gather_out_1_24 = 0;
localparam merge_in_1_24 = 1;
localparam gather_in_1_24 = 1;
localparam cast_sid_1_24 = 1022;
localparam gather_sid_1_24 = 0;

localparam cast_out_2_0 = 0;
localparam merge_out_2_0 = 0;
localparam gather_out_2_0 = 1;
localparam merge_in_2_0 = 0;
localparam gather_in_2_0 = 0;
localparam cast_sid_2_0 = 0;
localparam gather_sid_2_0 = 2;

localparam cast_out_2_1 = 1;
localparam merge_out_2_1 = 0;
localparam gather_out_2_1 = 0;
localparam merge_in_2_1 = 1;
localparam gather_in_2_1 = 0;
localparam cast_sid_2_1 = 15;
localparam gather_sid_2_1 = 0;

localparam cast_out_2_2 = 0;
localparam merge_out_2_2 = 1;
localparam gather_out_2_2 = 0;
localparam merge_in_2_2 = 0;
localparam gather_in_2_2 = 0;
localparam cast_sid_2_2 = 0;
localparam gather_sid_2_2 = 0;

localparam cast_out_2_3 = 0;
localparam merge_out_2_3 = 0;
localparam gather_out_2_3 = 1;
localparam merge_in_2_3 = 1;
localparam gather_in_2_3 = 0;
localparam cast_sid_2_3 = 0;
localparam gather_sid_2_3 = 17;

localparam cast_out_2_4 = 0;
localparam merge_out_2_4 = 1;
localparam gather_out_2_4 = 0;
localparam merge_in_2_4 = 0;
localparam gather_in_2_4 = 0;
localparam cast_sid_2_4 = 0;
localparam gather_sid_2_4 = 0;

localparam cast_out_2_5 = 1;
localparam merge_out_2_5 = 0;
localparam gather_out_2_5 = 1;
localparam merge_in_2_5 = 0;
localparam gather_in_2_5 = 1;
localparam cast_sid_2_5 = 38;
localparam gather_sid_2_5 = 23;

localparam cast_out_2_6 = 0;
localparam merge_out_2_6 = 1;
localparam gather_out_2_6 = 0;
localparam merge_in_2_6 = 0;
localparam gather_in_2_6 = 0;
localparam cast_sid_2_6 = 0;
localparam gather_sid_2_6 = 0;

localparam cast_out_2_7 = 1;
localparam merge_out_2_7 = 0;
localparam gather_out_2_7 = 1;
localparam merge_in_2_7 = 0;
localparam gather_in_2_7 = 1;
localparam cast_sid_2_7 = 50;
localparam gather_sid_2_7 = 31;

localparam cast_out_2_8 = 0;
localparam merge_out_2_8 = 1;
localparam gather_out_2_8 = 0;
localparam merge_in_2_8 = 0;
localparam gather_in_2_8 = 0;
localparam cast_sid_2_8 = 0;
localparam gather_sid_2_8 = 0;

localparam cast_out_2_9 = 1;
localparam merge_out_2_9 = 0;
localparam gather_out_2_9 = 0;
localparam merge_in_2_9 = 0;
localparam gather_in_2_9 = 1;
localparam cast_sid_2_9 = 62;
localparam gather_sid_2_9 = 0;

localparam cast_out_2_10 = 0;
localparam merge_out_2_10 = 1;
localparam gather_out_2_10 = 0;
localparam merge_in_2_10 = 0;
localparam gather_in_2_10 = 0;
localparam cast_sid_2_10 = 0;
localparam gather_sid_2_10 = 0;

localparam cast_out_2_11 = 0;
localparam merge_out_2_11 = 0;
localparam gather_out_2_11 = 1;
localparam merge_in_2_11 = 1;
localparam gather_in_2_11 = 0;
localparam cast_sid_2_11 = 0;
localparam gather_sid_2_11 = 46;

localparam cast_out_2_12 = 0;
localparam merge_out_2_12 = 1;
localparam gather_out_2_12 = 0;
localparam merge_in_2_12 = 0;
localparam gather_in_2_12 = 0;
localparam cast_sid_2_12 = 0;
localparam gather_sid_2_12 = 0;

localparam cast_out_2_13 = 0;
localparam merge_out_2_13 = 1;
localparam gather_out_2_13 = 0;
localparam merge_in_2_13 = 0;
localparam gather_in_2_13 = 0;
localparam cast_sid_2_13 = 0;
localparam gather_sid_2_13 = 0;

localparam cast_out_2_14 = 0;
localparam merge_out_2_14 = 1;
localparam gather_out_2_14 = 0;
localparam merge_in_2_14 = 0;
localparam gather_in_2_14 = 0;
localparam cast_sid_2_14 = 0;
localparam gather_sid_2_14 = 0;

localparam cast_out_2_15 = 0;
localparam merge_out_2_15 = 1;
localparam gather_out_2_15 = 0;
localparam merge_in_2_15 = 0;
localparam gather_in_2_15 = 0;
localparam cast_sid_2_15 = 0;
localparam gather_sid_2_15 = 0;

localparam cast_out_2_16 = 0;
localparam merge_out_2_16 = 1;
localparam gather_out_2_16 = 0;
localparam merge_in_2_16 = 0;
localparam gather_in_2_16 = 0;
localparam cast_sid_2_16 = 0;
localparam gather_sid_2_16 = 0;

localparam cast_out_2_17 = 0;
localparam merge_out_2_17 = 1;
localparam gather_out_2_17 = 0;
localparam merge_in_2_17 = 0;
localparam gather_in_2_17 = 0;
localparam cast_sid_2_17 = 0;
localparam gather_sid_2_17 = 0;

localparam cast_out_2_18 = 0;
localparam merge_out_2_18 = 1;
localparam gather_out_2_18 = 0;
localparam merge_in_2_18 = 0;
localparam gather_in_2_18 = 0;
localparam cast_sid_2_18 = 0;
localparam gather_sid_2_18 = 0;

localparam cast_out_2_19 = 0;
localparam merge_out_2_19 = 1;
localparam gather_out_2_19 = 0;
localparam merge_in_2_19 = 0;
localparam gather_in_2_19 = 0;
localparam cast_sid_2_19 = 0;
localparam gather_sid_2_19 = 0;

localparam cast_out_2_20 = 0;
localparam merge_out_2_20 = 1;
localparam gather_out_2_20 = 0;
localparam merge_in_2_20 = 0;
localparam gather_in_2_20 = 0;
localparam cast_sid_2_20 = 0;
localparam gather_sid_2_20 = 0;

localparam cast_out_2_21 = 0;
localparam merge_out_2_21 = 1;
localparam gather_out_2_21 = 0;
localparam merge_in_2_21 = 0;
localparam gather_in_2_21 = 0;
localparam cast_sid_2_21 = 0;
localparam gather_sid_2_21 = 0;

localparam cast_out_2_22 = 0;
localparam merge_out_2_22 = 1;
localparam gather_out_2_22 = 0;
localparam merge_in_2_22 = 0;
localparam gather_in_2_22 = 0;
localparam cast_sid_2_22 = 0;
localparam gather_sid_2_22 = 0;

localparam cast_out_2_23 = 0;
localparam merge_out_2_23 = 1;
localparam gather_out_2_23 = 0;
localparam merge_in_2_23 = 0;
localparam gather_in_2_23 = 0;
localparam cast_sid_2_23 = 0;
localparam gather_sid_2_23 = 0;

localparam cast_out_2_24 = 0;
localparam merge_out_2_24 = 0;
localparam gather_out_2_24 = 0;
localparam merge_in_2_24 = 0;
localparam gather_in_2_24 = 0;
localparam cast_sid_2_24 = 0;
localparam gather_sid_2_24 = 0;

localparam cast_out_3_0 = 1;
localparam merge_out_3_0 = 0;
localparam gather_out_3_0 = 0;
localparam merge_in_3_0 = 0;
localparam gather_in_3_0 = 0;
localparam cast_sid_3_0 = 3;
localparam gather_sid_3_0 = 0;

localparam cast_out_3_1 = 1;
localparam merge_out_3_1 = 0;
localparam gather_out_3_1 = 1;
localparam merge_in_3_1 = 0;
localparam gather_in_3_1 = 1;
localparam cast_sid_3_1 = 14;
localparam gather_sid_3_1 = 5;

localparam cast_out_3_2 = 1;
localparam merge_out_3_2 = 0;
localparam gather_out_3_2 = 0;
localparam merge_in_3_2 = 1;
localparam gather_in_3_2 = 0;
localparam cast_sid_3_2 = 19;
localparam gather_sid_3_2 = 0;

localparam cast_out_3_3 = 0;
localparam merge_out_3_3 = 1;
localparam gather_out_3_3 = 0;
localparam merge_in_3_3 = 0;
localparam gather_in_3_3 = 0;
localparam cast_sid_3_3 = 0;
localparam gather_sid_3_3 = 0;

localparam cast_out_3_4 = 1;
localparam merge_out_3_4 = 0;
localparam gather_out_3_4 = 0;
localparam merge_in_3_4 = 1;
localparam gather_in_3_4 = 0;
localparam cast_sid_3_4 = 28;
localparam gather_sid_3_4 = 0;

localparam cast_out_3_5 = 1;
localparam merge_out_3_5 = 0;
localparam gather_out_3_5 = 1;
localparam merge_in_3_5 = 0;
localparam gather_in_3_5 = 1;
localparam cast_sid_3_5 = 37;
localparam gather_sid_3_5 = 22;

localparam cast_out_3_6 = 1;
localparam merge_out_3_6 = 0;
localparam gather_out_3_6 = 0;
localparam merge_in_3_6 = 1;
localparam gather_in_3_6 = 0;
localparam cast_sid_3_6 = 40;
localparam gather_sid_3_6 = 0;

localparam cast_out_3_7 = 1;
localparam merge_out_3_7 = 0;
localparam gather_out_3_7 = 1;
localparam merge_in_3_7 = 0;
localparam gather_in_3_7 = 1;
localparam cast_sid_3_7 = 49;
localparam gather_sid_3_7 = 30;

localparam cast_out_3_8 = 1;
localparam merge_out_3_8 = 0;
localparam gather_out_3_8 = 0;
localparam merge_in_3_8 = 1;
localparam gather_in_3_8 = 0;
localparam cast_sid_3_8 = 52;
localparam gather_sid_3_8 = 0;

localparam cast_out_3_9 = 1;
localparam merge_out_3_9 = 0;
localparam gather_out_3_9 = 0;
localparam merge_in_3_9 = 0;
localparam gather_in_3_9 = 1;
localparam cast_sid_3_9 = 61;
localparam gather_sid_3_9 = 0;

localparam cast_out_3_10 = 0;
localparam merge_out_3_10 = 1;
localparam gather_out_3_10 = 0;
localparam merge_in_3_10 = 0;
localparam gather_in_3_10 = 0;
localparam cast_sid_3_10 = 0;
localparam gather_sid_3_10 = 0;

localparam cast_out_3_11 = 0;
localparam merge_out_3_11 = 1;
localparam gather_out_3_11 = 0;
localparam merge_in_3_11 = 0;
localparam gather_in_3_11 = 0;
localparam cast_sid_3_11 = 0;
localparam gather_sid_3_11 = 0;

localparam cast_out_3_12 = 0;
localparam merge_out_3_12 = 1;
localparam gather_out_3_12 = 0;
localparam merge_in_3_12 = 0;
localparam gather_in_3_12 = 0;
localparam cast_sid_3_12 = 0;
localparam gather_sid_3_12 = 0;

localparam cast_out_3_13 = 0;
localparam merge_out_3_13 = 0;
localparam gather_out_3_13 = 1;
localparam merge_in_3_13 = 1;
localparam gather_in_3_13 = 0;
localparam cast_sid_3_13 = 0;
localparam gather_sid_3_13 = 51;

localparam cast_out_3_14 = 0;
localparam merge_out_3_14 = 1;
localparam gather_out_3_14 = 0;
localparam merge_in_3_14 = 0;
localparam gather_in_3_14 = 0;
localparam cast_sid_3_14 = 0;
localparam gather_sid_3_14 = 0;

localparam cast_out_3_15 = 1;
localparam merge_out_3_15 = 0;
localparam gather_out_3_15 = 1;
localparam merge_in_3_15 = 1;
localparam gather_in_3_15 = 1;
localparam cast_sid_3_15 = 72;
localparam gather_sid_3_15 = 41;

localparam cast_out_3_16 = 0;
localparam merge_out_3_16 = 1;
localparam gather_out_3_16 = 0;
localparam merge_in_3_16 = 0;
localparam gather_in_3_16 = 0;
localparam cast_sid_3_16 = 0;
localparam gather_sid_3_16 = 0;

localparam cast_out_3_17 = 0;
localparam merge_out_3_17 = 1;
localparam gather_out_3_17 = 0;
localparam merge_in_3_17 = 0;
localparam gather_in_3_17 = 0;
localparam cast_sid_3_17 = 0;
localparam gather_sid_3_17 = 0;

localparam cast_out_3_18 = 0;
localparam merge_out_3_18 = 1;
localparam gather_out_3_18 = 0;
localparam merge_in_3_18 = 0;
localparam gather_in_3_18 = 0;
localparam cast_sid_3_18 = 0;
localparam gather_sid_3_18 = 0;

localparam cast_out_3_19 = 1;
localparam merge_out_3_19 = 0;
localparam gather_out_3_19 = 1;
localparam merge_in_3_19 = 1;
localparam gather_in_3_19 = 1;
localparam cast_sid_3_19 = 84;
localparam gather_sid_3_19 = 57;

localparam cast_out_3_20 = 0;
localparam merge_out_3_20 = 1;
localparam gather_out_3_20 = 0;
localparam merge_in_3_20 = 0;
localparam gather_in_3_20 = 0;
localparam cast_sid_3_20 = 0;
localparam gather_sid_3_20 = 0;

localparam cast_out_3_21 = 0;
localparam merge_out_3_21 = 1;
localparam gather_out_3_21 = 0;
localparam merge_in_3_21 = 0;
localparam gather_in_3_21 = 0;
localparam cast_sid_3_21 = 0;
localparam gather_sid_3_21 = 0;

localparam cast_out_3_22 = 0;
localparam merge_out_3_22 = 1;
localparam gather_out_3_22 = 0;
localparam merge_in_3_22 = 0;
localparam gather_in_3_22 = 0;
localparam cast_sid_3_22 = 0;
localparam gather_sid_3_22 = 0;

localparam cast_out_3_23 = 1;
localparam merge_out_3_23 = 0;
localparam gather_out_3_23 = 0;
localparam merge_in_3_23 = 1;
localparam gather_in_3_23 = 1;
localparam cast_sid_3_23 = 1022;
localparam gather_sid_3_23 = 0;

localparam cast_out_3_24 = 0;
localparam merge_out_3_24 = 0;
localparam gather_out_3_24 = 0;
localparam merge_in_3_24 = 0;
localparam gather_in_3_24 = 0;
localparam cast_sid_3_24 = 0;
localparam gather_sid_3_24 = 0;

localparam cast_out_4_0 = 1;
localparam merge_out_4_0 = 0;
localparam gather_out_4_0 = 1;
localparam merge_in_4_0 = 0;
localparam gather_in_4_0 = 1;
localparam cast_sid_4_0 = 4;
localparam gather_sid_4_0 = 1;

localparam cast_out_4_1 = 1;
localparam merge_out_4_1 = 0;
localparam gather_out_4_1 = 1;
localparam merge_in_4_1 = 0;
localparam gather_in_4_1 = 1;
localparam cast_sid_4_1 = 13;
localparam gather_sid_4_1 = 4;

localparam cast_out_4_2 = 1;
localparam merge_out_4_2 = 0;
localparam gather_out_4_2 = 0;
localparam merge_in_4_2 = 0;
localparam gather_in_4_2 = 0;
localparam cast_sid_4_2 = 20;
localparam gather_sid_4_2 = 0;

localparam cast_out_4_3 = 0;
localparam merge_out_4_3 = 0;
localparam gather_out_4_3 = 1;
localparam merge_in_4_3 = 1;
localparam gather_in_4_3 = 0;
localparam cast_sid_4_3 = 0;
localparam gather_sid_4_3 = 16;

localparam cast_out_4_4 = 1;
localparam merge_out_4_4 = 0;
localparam gather_out_4_4 = 1;
localparam merge_in_4_4 = 0;
localparam gather_in_4_4 = 1;
localparam cast_sid_4_4 = 29;
localparam gather_sid_4_4 = 12;

localparam cast_out_4_5 = 1;
localparam merge_out_4_5 = 0;
localparam gather_out_4_5 = 1;
localparam merge_in_4_5 = 0;
localparam gather_in_4_5 = 1;
localparam cast_sid_4_5 = 36;
localparam gather_sid_4_5 = 21;

localparam cast_out_4_6 = 1;
localparam merge_out_4_6 = 0;
localparam gather_out_4_6 = 1;
localparam merge_in_4_6 = 0;
localparam gather_in_4_6 = 1;
localparam cast_sid_4_6 = 41;
localparam gather_sid_4_6 = 24;

localparam cast_out_4_7 = 1;
localparam merge_out_4_7 = 0;
localparam gather_out_4_7 = 1;
localparam merge_in_4_7 = 0;
localparam gather_in_4_7 = 1;
localparam cast_sid_4_7 = 48;
localparam gather_sid_4_7 = 29;

localparam cast_out_4_8 = 1;
localparam merge_out_4_8 = 0;
localparam gather_out_4_8 = 1;
localparam merge_in_4_8 = 0;
localparam gather_in_4_8 = 1;
localparam cast_sid_4_8 = 53;
localparam gather_sid_4_8 = 32;

localparam cast_out_4_9 = 1;
localparam merge_out_4_9 = 0;
localparam gather_out_4_9 = 0;
localparam merge_in_4_9 = 0;
localparam gather_in_4_9 = 1;
localparam cast_sid_4_9 = 60;
localparam gather_sid_4_9 = 0;

localparam cast_out_4_10 = 0;
localparam merge_out_4_10 = 1;
localparam gather_out_4_10 = 0;
localparam merge_in_4_10 = 0;
localparam gather_in_4_10 = 0;
localparam cast_sid_4_10 = 0;
localparam gather_sid_4_10 = 0;

localparam cast_out_4_11 = 0;
localparam merge_out_4_11 = 1;
localparam gather_out_4_11 = 0;
localparam merge_in_4_11 = 0;
localparam gather_in_4_11 = 0;
localparam cast_sid_4_11 = 0;
localparam gather_sid_4_11 = 0;

localparam cast_out_4_12 = 0;
localparam merge_out_4_12 = 1;
localparam gather_out_4_12 = 0;
localparam merge_in_4_12 = 0;
localparam gather_in_4_12 = 0;
localparam cast_sid_4_12 = 0;
localparam gather_sid_4_12 = 0;

localparam cast_out_4_13 = 0;
localparam merge_out_4_13 = 1;
localparam gather_out_4_13 = 0;
localparam merge_in_4_13 = 0;
localparam gather_in_4_13 = 0;
localparam cast_sid_4_13 = 0;
localparam gather_sid_4_13 = 0;

localparam cast_out_4_14 = 0;
localparam merge_out_4_14 = 1;
localparam gather_out_4_14 = 0;
localparam merge_in_4_14 = 0;
localparam gather_in_4_14 = 0;
localparam cast_sid_4_14 = 0;
localparam gather_sid_4_14 = 0;

localparam cast_out_4_15 = 1;
localparam merge_out_4_15 = 0;
localparam gather_out_4_15 = 1;
localparam merge_in_4_15 = 1;
localparam gather_in_4_15 = 1;
localparam cast_sid_4_15 = 71;
localparam gather_sid_4_15 = 40;

localparam cast_out_4_16 = 0;
localparam merge_out_4_16 = 1;
localparam gather_out_4_16 = 0;
localparam merge_in_4_16 = 0;
localparam gather_in_4_16 = 0;
localparam cast_sid_4_16 = 0;
localparam gather_sid_4_16 = 0;

localparam cast_out_4_17 = 0;
localparam merge_out_4_17 = 1;
localparam gather_out_4_17 = 0;
localparam merge_in_4_17 = 0;
localparam gather_in_4_17 = 0;
localparam cast_sid_4_17 = 0;
localparam gather_sid_4_17 = 0;

localparam cast_out_4_18 = 0;
localparam merge_out_4_18 = 1;
localparam gather_out_4_18 = 0;
localparam merge_in_4_18 = 0;
localparam gather_in_4_18 = 0;
localparam cast_sid_4_18 = 0;
localparam gather_sid_4_18 = 0;

localparam cast_out_4_19 = 0;
localparam merge_out_4_19 = 1;
localparam gather_out_4_19 = 0;
localparam merge_in_4_19 = 0;
localparam gather_in_4_19 = 0;
localparam cast_sid_4_19 = 0;
localparam gather_sid_4_19 = 0;

localparam cast_out_4_20 = 0;
localparam merge_out_4_20 = 1;
localparam gather_out_4_20 = 0;
localparam merge_in_4_20 = 0;
localparam gather_in_4_20 = 0;
localparam cast_sid_4_20 = 0;
localparam gather_sid_4_20 = 0;

localparam cast_out_4_21 = 0;
localparam merge_out_4_21 = 1;
localparam gather_out_4_21 = 0;
localparam merge_in_4_21 = 0;
localparam gather_in_4_21 = 0;
localparam cast_sid_4_21 = 0;
localparam gather_sid_4_21 = 0;

localparam cast_out_4_22 = 0;
localparam merge_out_4_22 = 1;
localparam gather_out_4_22 = 0;
localparam merge_in_4_22 = 0;
localparam gather_in_4_22 = 0;
localparam cast_sid_4_22 = 0;
localparam gather_sid_4_22 = 0;

localparam cast_out_4_23 = 0;
localparam merge_out_4_23 = 1;
localparam gather_out_4_23 = 0;
localparam merge_in_4_23 = 0;
localparam gather_in_4_23 = 0;
localparam cast_sid_4_23 = 0;
localparam gather_sid_4_23 = 0;

localparam cast_out_4_24 = 0;
localparam merge_out_4_24 = 0;
localparam gather_out_4_24 = 0;
localparam merge_in_4_24 = 0;
localparam gather_in_4_24 = 0;
localparam cast_sid_4_24 = 0;
localparam gather_sid_4_24 = 0;

localparam cast_out_5_0 = 1;
localparam merge_out_5_0 = 0;
localparam gather_out_5_0 = 0;
localparam merge_in_5_0 = 0;
localparam gather_in_5_0 = 0;
localparam cast_sid_5_0 = 5;
localparam gather_sid_5_0 = 0;

localparam cast_out_5_1 = 1;
localparam merge_out_5_1 = 0;
localparam gather_out_5_1 = 0;
localparam merge_in_5_1 = 0;
localparam gather_in_5_1 = 0;
localparam cast_sid_5_1 = 12;
localparam gather_sid_5_1 = 0;

localparam cast_out_5_2 = 1;
localparam merge_out_5_2 = 0;
localparam gather_out_5_2 = 1;
localparam merge_in_5_2 = 0;
localparam gather_in_5_2 = 1;
localparam cast_sid_5_2 = 21;
localparam gather_sid_5_2 = 10;

localparam cast_out_5_3 = 0;
localparam merge_out_5_3 = 1;
localparam gather_out_5_3 = 0;
localparam merge_in_5_3 = 0;
localparam gather_in_5_3 = 0;
localparam cast_sid_5_3 = 0;
localparam gather_sid_5_3 = 0;

localparam cast_out_5_4 = 1;
localparam merge_out_5_4 = 0;
localparam gather_out_5_4 = 1;
localparam merge_in_5_4 = 0;
localparam gather_in_5_4 = 1;
localparam cast_sid_5_4 = 30;
localparam gather_sid_5_4 = 13;

localparam cast_out_5_5 = 1;
localparam merge_out_5_5 = 0;
localparam gather_out_5_5 = 1;
localparam merge_in_5_5 = 0;
localparam gather_in_5_5 = 1;
localparam cast_sid_5_5 = 35;
localparam gather_sid_5_5 = 20;

localparam cast_out_5_6 = 1;
localparam merge_out_5_6 = 0;
localparam gather_out_5_6 = 1;
localparam merge_in_5_6 = 0;
localparam gather_in_5_6 = 1;
localparam cast_sid_5_6 = 42;
localparam gather_sid_5_6 = 25;

localparam cast_out_5_7 = 1;
localparam merge_out_5_7 = 0;
localparam gather_out_5_7 = 1;
localparam merge_in_5_7 = 0;
localparam gather_in_5_7 = 1;
localparam cast_sid_5_7 = 47;
localparam gather_sid_5_7 = 28;

localparam cast_out_5_8 = 1;
localparam merge_out_5_8 = 0;
localparam gather_out_5_8 = 1;
localparam merge_in_5_8 = 0;
localparam gather_in_5_8 = 1;
localparam cast_sid_5_8 = 54;
localparam gather_sid_5_8 = 33;

localparam cast_out_5_9 = 1;
localparam merge_out_5_9 = 0;
localparam gather_out_5_9 = 0;
localparam merge_in_5_9 = 0;
localparam gather_in_5_9 = 1;
localparam cast_sid_5_9 = 59;
localparam gather_sid_5_9 = 0;

localparam cast_out_5_10 = 1;
localparam merge_out_5_10 = 0;
localparam gather_out_5_10 = 0;
localparam merge_in_5_10 = 1;
localparam gather_in_5_10 = 0;
localparam cast_sid_5_10 = 64;
localparam gather_sid_5_10 = 0;

localparam cast_out_5_11 = 0;
localparam merge_out_5_11 = 1;
localparam gather_out_5_11 = 0;
localparam merge_in_5_11 = 0;
localparam gather_in_5_11 = 0;
localparam cast_sid_5_11 = 0;
localparam gather_sid_5_11 = 0;

localparam cast_out_5_12 = 0;
localparam merge_out_5_12 = 0;
localparam gather_out_5_12 = 1;
localparam merge_in_5_12 = 1;
localparam gather_in_5_12 = 0;
localparam cast_sid_5_12 = 0;
localparam gather_sid_5_12 = 48;

localparam cast_out_5_13 = 0;
localparam merge_out_5_13 = 1;
localparam gather_out_5_13 = 0;
localparam merge_in_5_13 = 0;
localparam gather_in_5_13 = 0;
localparam cast_sid_5_13 = 0;
localparam gather_sid_5_13 = 0;

localparam cast_out_5_14 = 1;
localparam merge_out_5_14 = 0;
localparam gather_out_5_14 = 0;
localparam merge_in_5_14 = 1;
localparam gather_in_5_14 = 0;
localparam cast_sid_5_14 = 66;
localparam gather_sid_5_14 = 0;

localparam cast_out_5_15 = 0;
localparam merge_out_5_15 = 1;
localparam gather_out_5_15 = 0;
localparam merge_in_5_15 = 0;
localparam gather_in_5_15 = 0;
localparam cast_sid_5_15 = 0;
localparam gather_sid_5_15 = 0;

localparam cast_out_5_16 = 0;
localparam merge_out_5_16 = 1;
localparam gather_out_5_16 = 0;
localparam merge_in_5_16 = 0;
localparam gather_in_5_16 = 0;
localparam cast_sid_5_16 = 0;
localparam gather_sid_5_16 = 0;

localparam cast_out_5_17 = 0;
localparam merge_out_5_17 = 1;
localparam gather_out_5_17 = 0;
localparam merge_in_5_17 = 0;
localparam gather_in_5_17 = 0;
localparam cast_sid_5_17 = 0;
localparam gather_sid_5_17 = 0;

localparam cast_out_5_18 = 1;
localparam merge_out_5_18 = 0;
localparam gather_out_5_18 = 0;
localparam merge_in_5_18 = 1;
localparam gather_in_5_18 = 0;
localparam cast_sid_5_18 = 78;
localparam gather_sid_5_18 = 0;

localparam cast_out_5_19 = 1;
localparam merge_out_5_19 = 0;
localparam gather_out_5_19 = 1;
localparam merge_in_5_19 = 1;
localparam gather_in_5_19 = 1;
localparam cast_sid_5_19 = 83;
localparam gather_sid_5_19 = 56;

localparam cast_out_5_20 = 0;
localparam merge_out_5_20 = 1;
localparam gather_out_5_20 = 0;
localparam merge_in_5_20 = 0;
localparam gather_in_5_20 = 0;
localparam cast_sid_5_20 = 0;
localparam gather_sid_5_20 = 0;

localparam cast_out_5_21 = 1;
localparam merge_out_5_21 = 0;
localparam gather_out_5_21 = 0;
localparam merge_in_5_21 = 1;
localparam gather_in_5_21 = 0;
localparam cast_sid_5_21 = 88;
localparam gather_sid_5_21 = 0;

localparam cast_out_5_22 = 1;
localparam merge_out_5_22 = 0;
localparam gather_out_5_22 = 0;
localparam merge_in_5_22 = 1;
localparam gather_in_5_22 = 0;
localparam cast_sid_5_22 = 90;
localparam gather_sid_5_22 = 0;

localparam cast_out_5_23 = 1;
localparam merge_out_5_23 = 0;
localparam gather_out_5_23 = 0;
localparam merge_in_5_23 = 1;
localparam gather_in_5_23 = 1;
localparam cast_sid_5_23 = 1022;
localparam gather_sid_5_23 = 0;

localparam cast_out_5_24 = 0;
localparam merge_out_5_24 = 0;
localparam gather_out_5_24 = 0;
localparam merge_in_5_24 = 0;
localparam gather_in_5_24 = 0;
localparam cast_sid_5_24 = 0;
localparam gather_sid_5_24 = 0;

localparam cast_out_6_0 = 1;
localparam merge_out_6_0 = 0;
localparam gather_out_6_0 = 0;
localparam merge_in_6_0 = 0;
localparam gather_in_6_0 = 0;
localparam cast_sid_6_0 = 6;
localparam gather_sid_6_0 = 0;

localparam cast_out_6_1 = 0;
localparam merge_out_6_1 = 0;
localparam gather_out_6_1 = 1;
localparam merge_in_6_1 = 0;
localparam gather_in_6_1 = 0;
localparam cast_sid_6_1 = 0;
localparam gather_sid_6_1 = 7;

localparam cast_out_6_2 = 1;
localparam merge_out_6_2 = 0;
localparam gather_out_6_2 = 1;
localparam merge_in_6_2 = 0;
localparam gather_in_6_2 = 1;
localparam cast_sid_6_2 = 22;
localparam gather_sid_6_2 = 11;

localparam cast_out_6_3 = 1;
localparam merge_out_6_3 = 0;
localparam gather_out_6_3 = 0;
localparam merge_in_6_3 = 1;
localparam gather_in_6_3 = 0;
localparam cast_sid_6_3 = 27;
localparam gather_sid_6_3 = 0;

localparam cast_out_6_4 = 1;
localparam merge_out_6_4 = 0;
localparam gather_out_6_4 = 1;
localparam merge_in_6_4 = 0;
localparam gather_in_6_4 = 1;
localparam cast_sid_6_4 = 31;
localparam gather_sid_6_4 = 14;

localparam cast_out_6_5 = 1;
localparam merge_out_6_5 = 0;
localparam gather_out_6_5 = 0;
localparam merge_in_6_5 = 1;
localparam gather_in_6_5 = 0;
localparam cast_sid_6_5 = 34;
localparam gather_sid_6_5 = 0;

localparam cast_out_6_6 = 1;
localparam merge_out_6_6 = 0;
localparam gather_out_6_6 = 1;
localparam merge_in_6_6 = 0;
localparam gather_in_6_6 = 1;
localparam cast_sid_6_6 = 43;
localparam gather_sid_6_6 = 26;

localparam cast_out_6_7 = 0;
localparam merge_out_6_7 = 1;
localparam gather_out_6_7 = 0;
localparam merge_in_6_7 = 0;
localparam gather_in_6_7 = 0;
localparam cast_sid_6_7 = 0;
localparam gather_sid_6_7 = 0;

localparam cast_out_6_8 = 1;
localparam merge_out_6_8 = 0;
localparam gather_out_6_8 = 1;
localparam merge_in_6_8 = 0;
localparam gather_in_6_8 = 1;
localparam cast_sid_6_8 = 55;
localparam gather_sid_6_8 = 34;

localparam cast_out_6_9 = 1;
localparam merge_out_6_9 = 0;
localparam gather_out_6_9 = 0;
localparam merge_in_6_9 = 1;
localparam gather_in_6_9 = 0;
localparam cast_sid_6_9 = 58;
localparam gather_sid_6_9 = 0;

localparam cast_out_6_10 = 0;
localparam merge_out_6_10 = 1;
localparam gather_out_6_10 = 0;
localparam merge_in_6_10 = 0;
localparam gather_in_6_10 = 0;
localparam cast_sid_6_10 = 0;
localparam gather_sid_6_10 = 0;

localparam cast_out_6_11 = 0;
localparam merge_out_6_11 = 1;
localparam gather_out_6_11 = 0;
localparam merge_in_6_11 = 0;
localparam gather_in_6_11 = 0;
localparam cast_sid_6_11 = 0;
localparam gather_sid_6_11 = 0;

localparam cast_out_6_12 = 0;
localparam merge_out_6_12 = 1;
localparam gather_out_6_12 = 0;
localparam merge_in_6_12 = 0;
localparam gather_in_6_12 = 0;
localparam cast_sid_6_12 = 0;
localparam gather_sid_6_12 = 0;

localparam cast_out_6_13 = 0;
localparam merge_out_6_13 = 1;
localparam gather_out_6_13 = 0;
localparam merge_in_6_13 = 0;
localparam gather_in_6_13 = 0;
localparam cast_sid_6_13 = 0;
localparam gather_sid_6_13 = 0;

localparam cast_out_6_14 = 0;
localparam merge_out_6_14 = 1;
localparam gather_out_6_14 = 0;
localparam merge_in_6_14 = 0;
localparam gather_in_6_14 = 0;
localparam cast_sid_6_14 = 0;
localparam gather_sid_6_14 = 0;

localparam cast_out_6_15 = 1;
localparam merge_out_6_15 = 0;
localparam gather_out_6_15 = 1;
localparam merge_in_6_15 = 1;
localparam gather_in_6_15 = 1;
localparam cast_sid_6_15 = 70;
localparam gather_sid_6_15 = 39;

localparam cast_out_6_16 = 0;
localparam merge_out_6_16 = 1;
localparam gather_out_6_16 = 0;
localparam merge_in_6_16 = 0;
localparam gather_in_6_16 = 0;
localparam cast_sid_6_16 = 0;
localparam gather_sid_6_16 = 0;

localparam cast_out_6_17 = 1;
localparam merge_out_6_17 = 0;
localparam gather_out_6_17 = 0;
localparam merge_in_6_17 = 1;
localparam gather_in_6_17 = 0;
localparam cast_sid_6_17 = 76;
localparam gather_sid_6_17 = 0;

localparam cast_out_6_18 = 0;
localparam merge_out_6_18 = 1;
localparam gather_out_6_18 = 0;
localparam merge_in_6_18 = 0;
localparam gather_in_6_18 = 0;
localparam cast_sid_6_18 = 0;
localparam gather_sid_6_18 = 0;

localparam cast_out_6_19 = 1;
localparam merge_out_6_19 = 0;
localparam gather_out_6_19 = 1;
localparam merge_in_6_19 = 1;
localparam gather_in_6_19 = 1;
localparam cast_sid_6_19 = 82;
localparam gather_sid_6_19 = 55;

localparam cast_out_6_20 = 0;
localparam merge_out_6_20 = 1;
localparam gather_out_6_20 = 0;
localparam merge_in_6_20 = 0;
localparam gather_in_6_20 = 0;
localparam cast_sid_6_20 = 0;
localparam gather_sid_6_20 = 0;

localparam cast_out_6_21 = 0;
localparam merge_out_6_21 = 1;
localparam gather_out_6_21 = 0;
localparam merge_in_6_21 = 0;
localparam gather_in_6_21 = 0;
localparam cast_sid_6_21 = 0;
localparam gather_sid_6_21 = 0;

localparam cast_out_6_22 = 0;
localparam merge_out_6_22 = 1;
localparam gather_out_6_22 = 0;
localparam merge_in_6_22 = 0;
localparam gather_in_6_22 = 0;
localparam cast_sid_6_22 = 0;
localparam gather_sid_6_22 = 0;

localparam cast_out_6_23 = 1;
localparam merge_out_6_23 = 0;
localparam gather_out_6_23 = 0;
localparam merge_in_6_23 = 1;
localparam gather_in_6_23 = 1;
localparam cast_sid_6_23 = 1022;
localparam gather_sid_6_23 = 0;

localparam cast_out_6_24 = 0;
localparam merge_out_6_24 = 0;
localparam gather_out_6_24 = 0;
localparam merge_in_6_24 = 0;
localparam gather_in_6_24 = 0;
localparam cast_sid_6_24 = 0;
localparam gather_sid_6_24 = 0;

localparam cast_out_7_0 = 1;
localparam merge_out_7_0 = 0;
localparam gather_out_7_0 = 1;
localparam merge_in_7_0 = 0;
localparam gather_in_7_0 = 1;
localparam cast_sid_7_0 = 7;
localparam gather_sid_7_0 = 3;

localparam cast_out_7_1 = 0;
localparam merge_out_7_1 = 0;
localparam gather_out_7_1 = 1;
localparam merge_in_7_1 = 0;
localparam gather_in_7_1 = 0;
localparam cast_sid_7_1 = 0;
localparam gather_sid_7_1 = 6;

localparam cast_out_7_2 = 0;
localparam merge_out_7_2 = 1;
localparam gather_out_7_2 = 0;
localparam merge_in_7_2 = 0;
localparam gather_in_7_2 = 0;
localparam cast_sid_7_2 = 0;
localparam gather_sid_7_2 = 0;

localparam cast_out_7_3 = 0;
localparam merge_out_7_3 = 1;
localparam gather_out_7_3 = 0;
localparam merge_in_7_3 = 0;
localparam gather_in_7_3 = 0;
localparam cast_sid_7_3 = 0;
localparam gather_sid_7_3 = 0;

localparam cast_out_7_4 = 1;
localparam merge_out_7_4 = 0;
localparam gather_out_7_4 = 1;
localparam merge_in_7_4 = 0;
localparam gather_in_7_4 = 1;
localparam cast_sid_7_4 = 32;
localparam gather_sid_7_4 = 15;

localparam cast_out_7_5 = 0;
localparam merge_out_7_5 = 1;
localparam gather_out_7_5 = 0;
localparam merge_in_7_5 = 0;
localparam gather_in_7_5 = 0;
localparam cast_sid_7_5 = 0;
localparam gather_sid_7_5 = 0;

localparam cast_out_7_6 = 1;
localparam merge_out_7_6 = 0;
localparam gather_out_7_6 = 1;
localparam merge_in_7_6 = 0;
localparam gather_in_7_6 = 1;
localparam cast_sid_7_6 = 44;
localparam gather_sid_7_6 = 27;

localparam cast_out_7_7 = 1;
localparam merge_out_7_7 = 0;
localparam gather_out_7_7 = 0;
localparam merge_in_7_7 = 1;
localparam gather_in_7_7 = 0;
localparam cast_sid_7_7 = 46;
localparam gather_sid_7_7 = 0;

localparam cast_out_7_8 = 1;
localparam merge_out_7_8 = 0;
localparam gather_out_7_8 = 1;
localparam merge_in_7_8 = 0;
localparam gather_in_7_8 = 1;
localparam cast_sid_7_8 = 56;
localparam gather_sid_7_8 = 35;

localparam cast_out_7_9 = 0;
localparam merge_out_7_9 = 1;
localparam gather_out_7_9 = 0;
localparam merge_in_7_9 = 0;
localparam gather_in_7_9 = 0;
localparam cast_sid_7_9 = 0;
localparam gather_sid_7_9 = 0;

localparam cast_out_7_10 = 0;
localparam merge_out_7_10 = 1;
localparam gather_out_7_10 = 0;
localparam merge_in_7_10 = 0;
localparam gather_in_7_10 = 0;
localparam cast_sid_7_10 = 0;
localparam gather_sid_7_10 = 0;

localparam cast_out_7_11 = 0;
localparam merge_out_7_11 = 1;
localparam gather_out_7_11 = 0;
localparam merge_in_7_11 = 0;
localparam gather_in_7_11 = 0;
localparam cast_sid_7_11 = 0;
localparam gather_sid_7_11 = 0;

localparam cast_out_7_12 = 0;
localparam merge_out_7_12 = 1;
localparam gather_out_7_12 = 0;
localparam merge_in_7_12 = 0;
localparam gather_in_7_12 = 0;
localparam cast_sid_7_12 = 0;
localparam gather_sid_7_12 = 0;

localparam cast_out_7_13 = 0;
localparam merge_out_7_13 = 1;
localparam gather_out_7_13 = 0;
localparam merge_in_7_13 = 0;
localparam gather_in_7_13 = 0;
localparam cast_sid_7_13 = 0;
localparam gather_sid_7_13 = 0;

localparam cast_out_7_14 = 1;
localparam merge_out_7_14 = 0;
localparam gather_out_7_14 = 1;
localparam merge_in_7_14 = 1;
localparam gather_in_7_14 = 1;
localparam cast_sid_7_14 = 67;
localparam gather_sid_7_14 = 36;

localparam cast_out_7_15 = 0;
localparam merge_out_7_15 = 1;
localparam gather_out_7_15 = 0;
localparam merge_in_7_15 = 0;
localparam gather_in_7_15 = 0;
localparam cast_sid_7_15 = 0;
localparam gather_sid_7_15 = 0;

localparam cast_out_7_16 = 0;
localparam merge_out_7_16 = 1;
localparam gather_out_7_16 = 0;
localparam merge_in_7_16 = 0;
localparam gather_in_7_16 = 0;
localparam cast_sid_7_16 = 0;
localparam gather_sid_7_16 = 0;

localparam cast_out_7_17 = 0;
localparam merge_out_7_17 = 1;
localparam gather_out_7_17 = 0;
localparam merge_in_7_17 = 0;
localparam gather_in_7_17 = 0;
localparam cast_sid_7_17 = 0;
localparam gather_sid_7_17 = 0;

localparam cast_out_7_18 = 1;
localparam merge_out_7_18 = 0;
localparam gather_out_7_18 = 1;
localparam merge_in_7_18 = 1;
localparam gather_in_7_18 = 1;
localparam cast_sid_7_18 = 79;
localparam gather_sid_7_18 = 52;

localparam cast_out_7_19 = 0;
localparam merge_out_7_19 = 1;
localparam gather_out_7_19 = 0;
localparam merge_in_7_19 = 0;
localparam gather_in_7_19 = 0;
localparam cast_sid_7_19 = 0;
localparam gather_sid_7_19 = 0;

localparam cast_out_7_20 = 0;
localparam merge_out_7_20 = 1;
localparam gather_out_7_20 = 0;
localparam merge_in_7_20 = 0;
localparam gather_in_7_20 = 0;
localparam cast_sid_7_20 = 0;
localparam gather_sid_7_20 = 0;

localparam cast_out_7_21 = 0;
localparam merge_out_7_21 = 1;
localparam gather_out_7_21 = 0;
localparam merge_in_7_21 = 0;
localparam gather_in_7_21 = 0;
localparam cast_sid_7_21 = 0;
localparam gather_sid_7_21 = 0;

localparam cast_out_7_22 = 1;
localparam merge_out_7_22 = 0;
localparam gather_out_7_22 = 0;
localparam merge_in_7_22 = 1;
localparam gather_in_7_22 = 1;
localparam cast_sid_7_22 = 1022;
localparam gather_sid_7_22 = 0;

localparam cast_out_7_23 = 0;
localparam merge_out_7_23 = 1;
localparam gather_out_7_23 = 0;
localparam merge_in_7_23 = 0;
localparam gather_in_7_23 = 0;
localparam cast_sid_7_23 = 0;
localparam gather_sid_7_23 = 0;

localparam cast_out_7_24 = 0;
localparam merge_out_7_24 = 0;
localparam gather_out_7_24 = 0;
localparam merge_in_7_24 = 0;
localparam gather_in_7_24 = 0;
localparam cast_sid_7_24 = 0;
localparam gather_sid_7_24 = 0;

localparam cast_out_8_0 = 1;
localparam merge_out_8_0 = 0;
localparam gather_out_8_0 = 0;
localparam merge_in_8_0 = 0;
localparam gather_in_8_0 = 0;
localparam cast_sid_8_0 = 8;
localparam gather_sid_8_0 = 0;

localparam cast_out_8_1 = 1;
localparam merge_out_8_1 = 0;
localparam gather_out_8_1 = 0;
localparam merge_in_8_1 = 0;
localparam gather_in_8_1 = 0;
localparam cast_sid_8_1 = 11;
localparam gather_sid_8_1 = 0;

localparam cast_out_8_2 = 1;
localparam merge_out_8_2 = 0;
localparam gather_out_8_2 = 0;
localparam merge_in_8_2 = 1;
localparam gather_in_8_2 = 0;
localparam cast_sid_8_2 = 23;
localparam gather_sid_8_2 = 0;

localparam cast_out_8_3 = 1;
localparam merge_out_8_3 = 0;
localparam gather_out_8_3 = 0;
localparam merge_in_8_3 = 0;
localparam gather_in_8_3 = 1;
localparam cast_sid_8_3 = 26;
localparam gather_sid_8_3 = 0;

localparam cast_out_8_4 = 0;
localparam merge_out_8_4 = 1;
localparam gather_out_8_4 = 0;
localparam merge_in_8_4 = 0;
localparam gather_in_8_4 = 0;
localparam cast_sid_8_4 = 0;
localparam gather_sid_8_4 = 0;

localparam cast_out_8_5 = 1;
localparam merge_out_8_5 = 0;
localparam gather_out_8_5 = 0;
localparam merge_in_8_5 = 1;
localparam gather_in_8_5 = 0;
localparam cast_sid_8_5 = 33;
localparam gather_sid_8_5 = 0;

localparam cast_out_8_6 = 0;
localparam merge_out_8_6 = 1;
localparam gather_out_8_6 = 0;
localparam merge_in_8_6 = 0;
localparam gather_in_8_6 = 0;
localparam cast_sid_8_6 = 0;
localparam gather_sid_8_6 = 0;

localparam cast_out_8_7 = 0;
localparam merge_out_8_7 = 1;
localparam gather_out_8_7 = 0;
localparam merge_in_8_7 = 0;
localparam gather_in_8_7 = 0;
localparam cast_sid_8_7 = 0;
localparam gather_sid_8_7 = 0;

localparam cast_out_8_8 = 0;
localparam merge_out_8_8 = 1;
localparam gather_out_8_8 = 0;
localparam merge_in_8_8 = 0;
localparam gather_in_8_8 = 0;
localparam cast_sid_8_8 = 0;
localparam gather_sid_8_8 = 0;

localparam cast_out_8_9 = 0;
localparam merge_out_8_9 = 1;
localparam gather_out_8_9 = 0;
localparam merge_in_8_9 = 0;
localparam gather_in_8_9 = 0;
localparam cast_sid_8_9 = 0;
localparam gather_sid_8_9 = 0;

localparam cast_out_8_10 = 0;
localparam merge_out_8_10 = 1;
localparam gather_out_8_10 = 0;
localparam merge_in_8_10 = 0;
localparam gather_in_8_10 = 0;
localparam cast_sid_8_10 = 0;
localparam gather_sid_8_10 = 0;

localparam cast_out_8_11 = 0;
localparam merge_out_8_11 = 1;
localparam gather_out_8_11 = 0;
localparam merge_in_8_11 = 0;
localparam gather_in_8_11 = 0;
localparam cast_sid_8_11 = 0;
localparam gather_sid_8_11 = 0;

localparam cast_out_8_12 = 0;
localparam merge_out_8_12 = 1;
localparam gather_out_8_12 = 0;
localparam merge_in_8_12 = 0;
localparam gather_in_8_12 = 0;
localparam cast_sid_8_12 = 0;
localparam gather_sid_8_12 = 0;

localparam cast_out_8_13 = 0;
localparam merge_out_8_13 = 1;
localparam gather_out_8_13 = 0;
localparam merge_in_8_13 = 0;
localparam gather_in_8_13 = 0;
localparam cast_sid_8_13 = 0;
localparam gather_sid_8_13 = 0;

localparam cast_out_8_14 = 0;
localparam merge_out_8_14 = 1;
localparam gather_out_8_14 = 0;
localparam merge_in_8_14 = 0;
localparam gather_in_8_14 = 0;
localparam cast_sid_8_14 = 0;
localparam gather_sid_8_14 = 0;

localparam cast_out_8_15 = 1;
localparam merge_out_8_15 = 0;
localparam gather_out_8_15 = 1;
localparam merge_in_8_15 = 1;
localparam gather_in_8_15 = 1;
localparam cast_sid_8_15 = 69;
localparam gather_sid_8_15 = 38;

localparam cast_out_8_16 = 0;
localparam merge_out_8_16 = 1;
localparam gather_out_8_16 = 0;
localparam merge_in_8_16 = 0;
localparam gather_in_8_16 = 0;
localparam cast_sid_8_16 = 0;
localparam gather_sid_8_16 = 0;

localparam cast_out_8_17 = 0;
localparam merge_out_8_17 = 1;
localparam gather_out_8_17 = 0;
localparam merge_in_8_17 = 0;
localparam gather_in_8_17 = 0;
localparam cast_sid_8_17 = 0;
localparam gather_sid_8_17 = 0;

localparam cast_out_8_18 = 0;
localparam merge_out_8_18 = 1;
localparam gather_out_8_18 = 0;
localparam merge_in_8_18 = 0;
localparam gather_in_8_18 = 0;
localparam cast_sid_8_18 = 0;
localparam gather_sid_8_18 = 0;

localparam cast_out_8_19 = 0;
localparam merge_out_8_19 = 1;
localparam gather_out_8_19 = 0;
localparam merge_in_8_19 = 0;
localparam gather_in_8_19 = 0;
localparam cast_sid_8_19 = 0;
localparam gather_sid_8_19 = 0;

localparam cast_out_8_20 = 0;
localparam merge_out_8_20 = 1;
localparam gather_out_8_20 = 0;
localparam merge_in_8_20 = 0;
localparam gather_in_8_20 = 0;
localparam cast_sid_8_20 = 0;
localparam gather_sid_8_20 = 0;

localparam cast_out_8_21 = 0;
localparam merge_out_8_21 = 1;
localparam gather_out_8_21 = 0;
localparam merge_in_8_21 = 0;
localparam gather_in_8_21 = 0;
localparam cast_sid_8_21 = 0;
localparam gather_sid_8_21 = 0;

localparam cast_out_8_22 = 0;
localparam merge_out_8_22 = 1;
localparam gather_out_8_22 = 0;
localparam merge_in_8_22 = 0;
localparam gather_in_8_22 = 0;
localparam cast_sid_8_22 = 0;
localparam gather_sid_8_22 = 0;

localparam cast_out_8_23 = 1;
localparam merge_out_8_23 = 0;
localparam gather_out_8_23 = 0;
localparam merge_in_8_23 = 1;
localparam gather_in_8_23 = 1;
localparam cast_sid_8_23 = 1022;
localparam gather_sid_8_23 = 0;

localparam cast_out_8_24 = 0;
localparam merge_out_8_24 = 0;
localparam gather_out_8_24 = 0;
localparam merge_in_8_24 = 0;
localparam gather_in_8_24 = 0;
localparam cast_sid_8_24 = 0;
localparam gather_sid_8_24 = 0;

localparam cast_out_9_0 = 1;
localparam merge_out_9_0 = 0;
localparam gather_out_9_0 = 0;
localparam merge_in_9_0 = 0;
localparam gather_in_9_0 = 0;
localparam cast_sid_9_0 = 9;
localparam gather_sid_9_0 = 0;

localparam cast_out_9_1 = 1;
localparam merge_out_9_1 = 0;
localparam gather_out_9_1 = 0;
localparam merge_in_9_1 = 0;
localparam gather_in_9_1 = 1;
localparam cast_sid_9_1 = 10;
localparam gather_sid_9_1 = 0;

localparam cast_out_9_2 = 1;
localparam merge_out_9_2 = 0;
localparam gather_out_9_2 = 0;
localparam merge_in_9_2 = 0;
localparam gather_in_9_2 = 0;
localparam cast_sid_9_2 = 24;
localparam gather_sid_9_2 = 0;

localparam cast_out_9_3 = 1;
localparam merge_out_9_3 = 0;
localparam gather_out_9_3 = 0;
localparam merge_in_9_3 = 0;
localparam gather_in_9_3 = 1;
localparam cast_sid_9_3 = 25;
localparam gather_sid_9_3 = 0;

localparam cast_out_9_4 = 0;
localparam merge_out_9_4 = 1;
localparam gather_out_9_4 = 0;
localparam merge_in_9_4 = 0;
localparam gather_in_9_4 = 0;
localparam cast_sid_9_4 = 0;
localparam gather_sid_9_4 = 0;

localparam cast_out_9_5 = 0;
localparam merge_out_9_5 = 1;
localparam gather_out_9_5 = 0;
localparam merge_in_9_5 = 0;
localparam gather_in_9_5 = 0;
localparam cast_sid_9_5 = 0;
localparam gather_sid_9_5 = 0;

localparam cast_out_9_6 = 0;
localparam merge_out_9_6 = 1;
localparam gather_out_9_6 = 0;
localparam merge_in_9_6 = 0;
localparam gather_in_9_6 = 0;
localparam cast_sid_9_6 = 0;
localparam gather_sid_9_6 = 0;

localparam cast_out_9_7 = 1;
localparam merge_out_9_7 = 0;
localparam gather_out_9_7 = 0;
localparam merge_in_9_7 = 1;
localparam gather_in_9_7 = 0;
localparam cast_sid_9_7 = 45;
localparam gather_sid_9_7 = 0;

localparam cast_out_9_8 = 0;
localparam merge_out_9_8 = 1;
localparam gather_out_9_8 = 0;
localparam merge_in_9_8 = 0;
localparam gather_in_9_8 = 0;
localparam cast_sid_9_8 = 0;
localparam gather_sid_9_8 = 0;

localparam cast_out_9_9 = 1;
localparam merge_out_9_9 = 0;
localparam gather_out_9_9 = 0;
localparam merge_in_9_9 = 1;
localparam gather_in_9_9 = 0;
localparam cast_sid_9_9 = 57;
localparam gather_sid_9_9 = 0;

localparam cast_out_9_10 = 0;
localparam merge_out_9_10 = 0;
localparam gather_out_9_10 = 1;
localparam merge_in_9_10 = 1;
localparam gather_in_9_10 = 0;
localparam cast_sid_9_10 = 0;
localparam gather_sid_9_10 = 44;

localparam cast_out_9_11 = 0;
localparam merge_out_9_11 = 0;
localparam gather_out_9_11 = 1;
localparam merge_in_9_11 = 1;
localparam gather_in_9_11 = 0;
localparam cast_sid_9_11 = 0;
localparam gather_sid_9_11 = 45;

localparam cast_out_9_12 = 0;
localparam merge_out_9_12 = 0;
localparam gather_out_9_12 = 1;
localparam merge_in_9_12 = 1;
localparam gather_in_9_12 = 0;
localparam cast_sid_9_12 = 0;
localparam gather_sid_9_12 = 49;

localparam cast_out_9_13 = 0;
localparam merge_out_9_13 = 0;
localparam gather_out_9_13 = 1;
localparam merge_in_9_13 = 1;
localparam gather_in_9_13 = 0;
localparam cast_sid_9_13 = 0;
localparam gather_sid_9_13 = 50;

localparam cast_out_9_14 = 1;
localparam merge_out_9_14 = 0;
localparam gather_out_9_14 = 1;
localparam merge_in_9_14 = 1;
localparam gather_in_9_14 = 1;
localparam cast_sid_9_14 = 68;
localparam gather_sid_9_14 = 37;

localparam cast_out_9_15 = 0;
localparam merge_out_9_15 = 1;
localparam gather_out_9_15 = 0;
localparam merge_in_9_15 = 0;
localparam gather_in_9_15 = 0;
localparam cast_sid_9_15 = 0;
localparam gather_sid_9_15 = 0;

localparam cast_out_9_16 = 1;
localparam merge_out_9_16 = 0;
localparam gather_out_9_16 = 0;
localparam merge_in_9_16 = 1;
localparam gather_in_9_16 = 0;
localparam cast_sid_9_16 = 75;
localparam gather_sid_9_16 = 0;

localparam cast_out_9_17 = 0;
localparam merge_out_9_17 = 1;
localparam gather_out_9_17 = 0;
localparam merge_in_9_17 = 0;
localparam gather_in_9_17 = 0;
localparam cast_sid_9_17 = 0;
localparam gather_sid_9_17 = 0;

localparam cast_out_9_18 = 1;
localparam merge_out_9_18 = 0;
localparam gather_out_9_18 = 1;
localparam merge_in_9_18 = 1;
localparam gather_in_9_18 = 1;
localparam cast_sid_9_18 = 80;
localparam gather_sid_9_18 = 53;

localparam cast_out_9_19 = 1;
localparam merge_out_9_19 = 0;
localparam gather_out_9_19 = 1;
localparam merge_in_9_19 = 1;
localparam gather_in_9_19 = 1;
localparam cast_sid_9_19 = 81;
localparam gather_sid_9_19 = 54;

localparam cast_out_9_20 = 1;
localparam merge_out_9_20 = 0;
localparam gather_out_9_20 = 0;
localparam merge_in_9_20 = 1;
localparam gather_in_9_20 = 0;
localparam cast_sid_9_20 = 87;
localparam gather_sid_9_20 = 0;

localparam cast_out_9_21 = 0;
localparam merge_out_9_21 = 1;
localparam gather_out_9_21 = 0;
localparam merge_in_9_21 = 0;
localparam gather_in_9_21 = 0;
localparam cast_sid_9_21 = 0;
localparam gather_sid_9_21 = 0;

localparam cast_out_9_22 = 1;
localparam merge_out_9_22 = 0;
localparam gather_out_9_22 = 0;
localparam merge_in_9_22 = 1;
localparam gather_in_9_22 = 1;
localparam cast_sid_9_22 = 1022;
localparam gather_sid_9_22 = 0;

localparam cast_out_9_23 = 0;
localparam merge_out_9_23 = 1;
localparam gather_out_9_23 = 0;
localparam merge_in_9_23 = 0;
localparam gather_in_9_23 = 0;
localparam cast_sid_9_23 = 0;
localparam gather_sid_9_23 = 0;

localparam cast_out_9_24 = 0;
localparam merge_out_9_24 = 0;
localparam gather_out_9_24 = 0;
localparam merge_in_9_24 = 0;
localparam gather_in_9_24 = 0;
localparam cast_sid_9_24 = 0;
localparam gather_sid_9_24 = 0;

`endif

