
//Merge Network
//Width: 5
//Height:6
`include "params.svh"
`include "merge_config.svh"

module merge_network(
    input       wire                            clk,
    input       wire                            rstn,

    //router local ports
    input       wire        [`DW-1:0]           data_i[`NOC_WIDTH][`NOC_HEIGHT],
    input       wire                            valid_i[`NOC_WIDTH][`NOC_HEIGHT],
    output      reg                             ready_o[`NOC_WIDTH][`NOC_HEIGHT],

    output      reg         [`DW-1:0]           data_o[`NOC_WIDTH][`NOC_HEIGHT],
    output      reg                             valid_o[`NOC_WIDTH][`NOC_HEIGHT],
    input       wire                            ready_i[`NOC_WIDTH][`NOC_HEIGHT]
);

reg [`DW-1:0] data_i_0_0[5];
reg valid_i_0_0[5], ready_i_0_0[5];    
wire [`DW-1:0] data_o_0_0[5];
wire valid_o_0_0[5], ready_o_0_0[5];        

reg [`DW-1:0] data_i_0_1[5];
reg valid_i_0_1[5], ready_i_0_1[5];    
wire [`DW-1:0] data_o_0_1[5];
wire valid_o_0_1[5], ready_o_0_1[5];        

reg [`DW-1:0] data_i_0_2[5];
reg valid_i_0_2[5], ready_i_0_2[5];    
wire [`DW-1:0] data_o_0_2[5];
wire valid_o_0_2[5], ready_o_0_2[5];        

reg [`DW-1:0] data_i_0_3[5];
reg valid_i_0_3[5], ready_i_0_3[5];    
wire [`DW-1:0] data_o_0_3[5];
wire valid_o_0_3[5], ready_o_0_3[5];        

reg [`DW-1:0] data_i_0_4[5];
reg valid_i_0_4[5], ready_i_0_4[5];    
wire [`DW-1:0] data_o_0_4[5];
wire valid_o_0_4[5], ready_o_0_4[5];        

reg [`DW-1:0] data_i_0_5[5];
reg valid_i_0_5[5], ready_i_0_5[5];    
wire [`DW-1:0] data_o_0_5[5];
wire valid_o_0_5[5], ready_o_0_5[5];        

reg [`DW-1:0] data_i_1_0[5];
reg valid_i_1_0[5], ready_i_1_0[5];    
wire [`DW-1:0] data_o_1_0[5];
wire valid_o_1_0[5], ready_o_1_0[5];        

reg [`DW-1:0] data_i_1_1[5];
reg valid_i_1_1[5], ready_i_1_1[5];    
wire [`DW-1:0] data_o_1_1[5];
wire valid_o_1_1[5], ready_o_1_1[5];        

reg [`DW-1:0] data_i_1_2[5];
reg valid_i_1_2[5], ready_i_1_2[5];    
wire [`DW-1:0] data_o_1_2[5];
wire valid_o_1_2[5], ready_o_1_2[5];        

reg [`DW-1:0] data_i_1_3[5];
reg valid_i_1_3[5], ready_i_1_3[5];    
wire [`DW-1:0] data_o_1_3[5];
wire valid_o_1_3[5], ready_o_1_3[5];        

reg [`DW-1:0] data_i_1_4[5];
reg valid_i_1_4[5], ready_i_1_4[5];    
wire [`DW-1:0] data_o_1_4[5];
wire valid_o_1_4[5], ready_o_1_4[5];        

reg [`DW-1:0] data_i_1_5[5];
reg valid_i_1_5[5], ready_i_1_5[5];    
wire [`DW-1:0] data_o_1_5[5];
wire valid_o_1_5[5], ready_o_1_5[5];        

reg [`DW-1:0] data_i_2_0[5];
reg valid_i_2_0[5], ready_i_2_0[5];    
wire [`DW-1:0] data_o_2_0[5];
wire valid_o_2_0[5], ready_o_2_0[5];        

reg [`DW-1:0] data_i_2_1[5];
reg valid_i_2_1[5], ready_i_2_1[5];    
wire [`DW-1:0] data_o_2_1[5];
wire valid_o_2_1[5], ready_o_2_1[5];        

reg [`DW-1:0] data_i_2_2[5];
reg valid_i_2_2[5], ready_i_2_2[5];    
wire [`DW-1:0] data_o_2_2[5];
wire valid_o_2_2[5], ready_o_2_2[5];        

reg [`DW-1:0] data_i_2_3[5];
reg valid_i_2_3[5], ready_i_2_3[5];    
wire [`DW-1:0] data_o_2_3[5];
wire valid_o_2_3[5], ready_o_2_3[5];        

reg [`DW-1:0] data_i_2_4[5];
reg valid_i_2_4[5], ready_i_2_4[5];    
wire [`DW-1:0] data_o_2_4[5];
wire valid_o_2_4[5], ready_o_2_4[5];        

reg [`DW-1:0] data_i_2_5[5];
reg valid_i_2_5[5], ready_i_2_5[5];    
wire [`DW-1:0] data_o_2_5[5];
wire valid_o_2_5[5], ready_o_2_5[5];        

reg [`DW-1:0] data_i_3_0[5];
reg valid_i_3_0[5], ready_i_3_0[5];    
wire [`DW-1:0] data_o_3_0[5];
wire valid_o_3_0[5], ready_o_3_0[5];        

reg [`DW-1:0] data_i_3_1[5];
reg valid_i_3_1[5], ready_i_3_1[5];    
wire [`DW-1:0] data_o_3_1[5];
wire valid_o_3_1[5], ready_o_3_1[5];        

reg [`DW-1:0] data_i_3_2[5];
reg valid_i_3_2[5], ready_i_3_2[5];    
wire [`DW-1:0] data_o_3_2[5];
wire valid_o_3_2[5], ready_o_3_2[5];        

reg [`DW-1:0] data_i_3_3[5];
reg valid_i_3_3[5], ready_i_3_3[5];    
wire [`DW-1:0] data_o_3_3[5];
wire valid_o_3_3[5], ready_o_3_3[5];        

reg [`DW-1:0] data_i_3_4[5];
reg valid_i_3_4[5], ready_i_3_4[5];    
wire [`DW-1:0] data_o_3_4[5];
wire valid_o_3_4[5], ready_o_3_4[5];        

reg [`DW-1:0] data_i_3_5[5];
reg valid_i_3_5[5], ready_i_3_5[5];    
wire [`DW-1:0] data_o_3_5[5];
wire valid_o_3_5[5], ready_o_3_5[5];        

reg [`DW-1:0] data_i_4_0[5];
reg valid_i_4_0[5], ready_i_4_0[5];    
wire [`DW-1:0] data_o_4_0[5];
wire valid_o_4_0[5], ready_o_4_0[5];        

reg [`DW-1:0] data_i_4_1[5];
reg valid_i_4_1[5], ready_i_4_1[5];    
wire [`DW-1:0] data_o_4_1[5];
wire valid_o_4_1[5], ready_o_4_1[5];        

reg [`DW-1:0] data_i_4_2[5];
reg valid_i_4_2[5], ready_i_4_2[5];    
wire [`DW-1:0] data_o_4_2[5];
wire valid_o_4_2[5], ready_o_4_2[5];        

reg [`DW-1:0] data_i_4_3[5];
reg valid_i_4_3[5], ready_i_4_3[5];    
wire [`DW-1:0] data_o_4_3[5];
wire valid_o_4_3[5], ready_o_4_3[5];        

reg [`DW-1:0] data_i_4_4[5];
reg valid_i_4_4[5], ready_i_4_4[5];    
wire [`DW-1:0] data_o_4_4[5];
wire valid_o_4_4[5], ready_o_4_4[5];        

reg [`DW-1:0] data_i_4_5[5];
reg valid_i_4_5[5], ready_i_4_5[5];    
wire [`DW-1:0] data_o_4_5[5];
wire valid_o_4_5[5], ready_o_4_5[5];        

always@(*) begin
    data_o[0][0] = data_o_0_0[0];
    valid_o[0][0] = valid_o_0_0[0];
    ready_o[0][0] = ready_o_0_0[0];
    data_o[0][1] = data_o_0_1[0];
    valid_o[0][1] = valid_o_0_1[0];
    ready_o[0][1] = ready_o_0_1[0];
    data_o[0][2] = data_o_0_2[0];
    valid_o[0][2] = valid_o_0_2[0];
    ready_o[0][2] = ready_o_0_2[0];
    data_o[0][3] = data_o_0_3[0];
    valid_o[0][3] = valid_o_0_3[0];
    ready_o[0][3] = ready_o_0_3[0];
    data_o[0][4] = data_o_0_4[0];
    valid_o[0][4] = valid_o_0_4[0];
    ready_o[0][4] = ready_o_0_4[0];
    data_o[0][5] = data_o_0_5[0];
    valid_o[0][5] = valid_o_0_5[0];
    ready_o[0][5] = ready_o_0_5[0];
    data_o[1][0] = data_o_1_0[0];
    valid_o[1][0] = valid_o_1_0[0];
    ready_o[1][0] = ready_o_1_0[0];
    data_o[1][1] = data_o_1_1[0];
    valid_o[1][1] = valid_o_1_1[0];
    ready_o[1][1] = ready_o_1_1[0];
    data_o[1][2] = data_o_1_2[0];
    valid_o[1][2] = valid_o_1_2[0];
    ready_o[1][2] = ready_o_1_2[0];
    data_o[1][3] = data_o_1_3[0];
    valid_o[1][3] = valid_o_1_3[0];
    ready_o[1][3] = ready_o_1_3[0];
    data_o[1][4] = data_o_1_4[0];
    valid_o[1][4] = valid_o_1_4[0];
    ready_o[1][4] = ready_o_1_4[0];
    data_o[1][5] = data_o_1_5[0];
    valid_o[1][5] = valid_o_1_5[0];
    ready_o[1][5] = ready_o_1_5[0];
    data_o[2][0] = data_o_2_0[0];
    valid_o[2][0] = valid_o_2_0[0];
    ready_o[2][0] = ready_o_2_0[0];
    data_o[2][1] = data_o_2_1[0];
    valid_o[2][1] = valid_o_2_1[0];
    ready_o[2][1] = ready_o_2_1[0];
    data_o[2][2] = data_o_2_2[0];
    valid_o[2][2] = valid_o_2_2[0];
    ready_o[2][2] = ready_o_2_2[0];
    data_o[2][3] = data_o_2_3[0];
    valid_o[2][3] = valid_o_2_3[0];
    ready_o[2][3] = ready_o_2_3[0];
    data_o[2][4] = data_o_2_4[0];
    valid_o[2][4] = valid_o_2_4[0];
    ready_o[2][4] = ready_o_2_4[0];
    data_o[2][5] = data_o_2_5[0];
    valid_o[2][5] = valid_o_2_5[0];
    ready_o[2][5] = ready_o_2_5[0];
    data_o[3][0] = data_o_3_0[0];
    valid_o[3][0] = valid_o_3_0[0];
    ready_o[3][0] = ready_o_3_0[0];
    data_o[3][1] = data_o_3_1[0];
    valid_o[3][1] = valid_o_3_1[0];
    ready_o[3][1] = ready_o_3_1[0];
    data_o[3][2] = data_o_3_2[0];
    valid_o[3][2] = valid_o_3_2[0];
    ready_o[3][2] = ready_o_3_2[0];
    data_o[3][3] = data_o_3_3[0];
    valid_o[3][3] = valid_o_3_3[0];
    ready_o[3][3] = ready_o_3_3[0];
    data_o[3][4] = data_o_3_4[0];
    valid_o[3][4] = valid_o_3_4[0];
    ready_o[3][4] = ready_o_3_4[0];
    data_o[3][5] = data_o_3_5[0];
    valid_o[3][5] = valid_o_3_5[0];
    ready_o[3][5] = ready_o_3_5[0];
    data_o[4][0] = data_o_4_0[0];
    valid_o[4][0] = valid_o_4_0[0];
    ready_o[4][0] = ready_o_4_0[0];
    data_o[4][1] = data_o_4_1[0];
    valid_o[4][1] = valid_o_4_1[0];
    ready_o[4][1] = ready_o_4_1[0];
    data_o[4][2] = data_o_4_2[0];
    valid_o[4][2] = valid_o_4_2[0];
    ready_o[4][2] = ready_o_4_2[0];
    data_o[4][3] = data_o_4_3[0];
    valid_o[4][3] = valid_o_4_3[0];
    ready_o[4][3] = ready_o_4_3[0];
    data_o[4][4] = data_o_4_4[0];
    valid_o[4][4] = valid_o_4_4[0];
    ready_o[4][4] = ready_o_4_4[0];
    data_o[4][5] = data_o_4_5[0];
    valid_o[4][5] = valid_o_4_5[0];
    ready_o[4][5] = ready_o_4_5[0];
end

/*Router 0,0*/    
merge_router #(
    .input_mask                     (input_mask_0_0),
    .output_sel                     (output_sel_0_0)
)router0(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_0_0),
    .valid_i                        (valid_i_0_0),
    .ready_o                        (ready_o_0_0),
    .data_o                         (data_o_0_0),
    .valid_o                        (valid_o_0_0),
    .ready_i                        (ready_i_0_0)
);


always@(*) begin
    data_i_0_0[4] = data_o_0_1[3];
    valid_i_0_0[4] = valid_o_0_1[3];
    ready_i_0_0[4] = ready_o_0_1[3];
    data_i_0_0[2] = data_o_1_0[1];
    valid_i_0_0[2] = valid_o_1_0[1];
    ready_i_0_0[2] = ready_o_1_0[1];
    data_i_0_0[0] = data_i[0][0];
    valid_i_0_0[0] = valid_i[0][0];
    ready_i_0_0[0] = ready_i[0][0];
end


/*Router 0,1*/    
merge_router #(
    .input_mask                     (input_mask_0_1),
    .output_sel                     (output_sel_0_1)
)router5(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_0_1),
    .valid_i                        (valid_i_0_1),
    .ready_o                        (ready_o_0_1),
    .data_o                         (data_o_0_1),
    .valid_o                        (valid_o_0_1),
    .ready_i                        (ready_i_0_1)
);


always@(*) begin
    data_i_0_1[3] = data_o_0_0[4];
    valid_i_0_1[3] = valid_o_0_0[4];
    ready_i_0_1[3] = ready_o_0_0[4];
    data_i_0_1[4] = data_o_0_2[3];
    valid_i_0_1[4] = valid_o_0_2[3];
    ready_i_0_1[4] = ready_o_0_2[3];
    data_i_0_1[2] = data_o_1_1[1];
    valid_i_0_1[2] = valid_o_1_1[1];
    ready_i_0_1[2] = ready_o_1_1[1];
    data_i_0_1[0] = data_i[0][1];
    valid_i_0_1[0] = valid_i[0][1];
    ready_i_0_1[0] = ready_i[0][1];
end


/*Router 0,2*/    
merge_router #(
    .input_mask                     (input_mask_0_2),
    .output_sel                     (output_sel_0_2)
)router10(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_0_2),
    .valid_i                        (valid_i_0_2),
    .ready_o                        (ready_o_0_2),
    .data_o                         (data_o_0_2),
    .valid_o                        (valid_o_0_2),
    .ready_i                        (ready_i_0_2)
);


always@(*) begin
    data_i_0_2[3] = data_o_0_1[4];
    valid_i_0_2[3] = valid_o_0_1[4];
    ready_i_0_2[3] = ready_o_0_1[4];
    data_i_0_2[4] = data_o_0_3[3];
    valid_i_0_2[4] = valid_o_0_3[3];
    ready_i_0_2[4] = ready_o_0_3[3];
    data_i_0_2[2] = data_o_1_2[1];
    valid_i_0_2[2] = valid_o_1_2[1];
    ready_i_0_2[2] = ready_o_1_2[1];
    data_i_0_2[0] = data_i[0][2];
    valid_i_0_2[0] = valid_i[0][2];
    ready_i_0_2[0] = ready_i[0][2];
end


/*Router 0,3*/    
merge_router #(
    .input_mask                     (input_mask_0_3),
    .output_sel                     (output_sel_0_3)
)router15(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_0_3),
    .valid_i                        (valid_i_0_3),
    .ready_o                        (ready_o_0_3),
    .data_o                         (data_o_0_3),
    .valid_o                        (valid_o_0_3),
    .ready_i                        (ready_i_0_3)
);


always@(*) begin
    data_i_0_3[3] = data_o_0_2[4];
    valid_i_0_3[3] = valid_o_0_2[4];
    ready_i_0_3[3] = ready_o_0_2[4];
    data_i_0_3[4] = data_o_0_4[3];
    valid_i_0_3[4] = valid_o_0_4[3];
    ready_i_0_3[4] = ready_o_0_4[3];
    data_i_0_3[2] = data_o_1_3[1];
    valid_i_0_3[2] = valid_o_1_3[1];
    ready_i_0_3[2] = ready_o_1_3[1];
    data_i_0_3[0] = data_i[0][3];
    valid_i_0_3[0] = valid_i[0][3];
    ready_i_0_3[0] = ready_i[0][3];
end


/*Router 0,4*/    
merge_router #(
    .input_mask                     (input_mask_0_4),
    .output_sel                     (output_sel_0_4)
)router20(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_0_4),
    .valid_i                        (valid_i_0_4),
    .ready_o                        (ready_o_0_4),
    .data_o                         (data_o_0_4),
    .valid_o                        (valid_o_0_4),
    .ready_i                        (ready_i_0_4)
);


always@(*) begin
    data_i_0_4[3] = data_o_0_3[4];
    valid_i_0_4[3] = valid_o_0_3[4];
    ready_i_0_4[3] = ready_o_0_3[4];
    data_i_0_4[4] = data_o_0_5[3];
    valid_i_0_4[4] = valid_o_0_5[3];
    ready_i_0_4[4] = ready_o_0_5[3];
    data_i_0_4[2] = data_o_1_4[1];
    valid_i_0_4[2] = valid_o_1_4[1];
    ready_i_0_4[2] = ready_o_1_4[1];
    data_i_0_4[0] = data_i[0][4];
    valid_i_0_4[0] = valid_i[0][4];
    ready_i_0_4[0] = ready_i[0][4];
end


/*Router 0,5*/    
merge_router #(
    .input_mask                     (input_mask_0_5),
    .output_sel                     (output_sel_0_5)
)router25(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_0_5),
    .valid_i                        (valid_i_0_5),
    .ready_o                        (ready_o_0_5),
    .data_o                         (data_o_0_5),
    .valid_o                        (valid_o_0_5),
    .ready_i                        (ready_i_0_5)
);


always@(*) begin
    data_i_0_5[3] = data_o_0_4[4];
    valid_i_0_5[3] = valid_o_0_4[4];
    ready_i_0_5[3] = ready_o_0_4[4];
    data_i_0_5[2] = data_o_1_5[1];
    valid_i_0_5[2] = valid_o_1_5[1];
    ready_i_0_5[2] = ready_o_1_5[1];
    data_i_0_5[0] = data_i[0][5];
    valid_i_0_5[0] = valid_i[0][5];
    ready_i_0_5[0] = ready_i[0][5];
end


/*Router 1,0*/    
merge_router #(
    .input_mask                     (input_mask_1_0),
    .output_sel                     (output_sel_1_0)
)router1(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_1_0),
    .valid_i                        (valid_i_1_0),
    .ready_o                        (ready_o_1_0),
    .data_o                         (data_o_1_0),
    .valid_o                        (valid_o_1_0),
    .ready_i                        (ready_i_1_0)
);


always@(*) begin
    data_i_1_0[4] = data_o_1_1[3];
    valid_i_1_0[4] = valid_o_1_1[3];
    ready_i_1_0[4] = ready_o_1_1[3];
    data_i_1_0[1] = data_o_0_0[2];
    valid_i_1_0[1] = valid_o_0_0[2];
    ready_i_1_0[1] = ready_o_0_0[2];
    data_i_1_0[2] = data_o_2_0[1];
    valid_i_1_0[2] = valid_o_2_0[1];
    ready_i_1_0[2] = ready_o_2_0[1];
    data_i_1_0[0] = data_i[1][0];
    valid_i_1_0[0] = valid_i[1][0];
    ready_i_1_0[0] = ready_i[1][0];
end


/*Router 1,1*/    
merge_router #(
    .input_mask                     (input_mask_1_1),
    .output_sel                     (output_sel_1_1)
)router6(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_1_1),
    .valid_i                        (valid_i_1_1),
    .ready_o                        (ready_o_1_1),
    .data_o                         (data_o_1_1),
    .valid_o                        (valid_o_1_1),
    .ready_i                        (ready_i_1_1)
);


always@(*) begin
    data_i_1_1[3] = data_o_1_0[4];
    valid_i_1_1[3] = valid_o_1_0[4];
    ready_i_1_1[3] = ready_o_1_0[4];
    data_i_1_1[4] = data_o_1_2[3];
    valid_i_1_1[4] = valid_o_1_2[3];
    ready_i_1_1[4] = ready_o_1_2[3];
    data_i_1_1[1] = data_o_0_1[2];
    valid_i_1_1[1] = valid_o_0_1[2];
    ready_i_1_1[1] = ready_o_0_1[2];
    data_i_1_1[2] = data_o_2_1[1];
    valid_i_1_1[2] = valid_o_2_1[1];
    ready_i_1_1[2] = ready_o_2_1[1];
    data_i_1_1[0] = data_i[1][1];
    valid_i_1_1[0] = valid_i[1][1];
    ready_i_1_1[0] = ready_i[1][1];
end


/*Router 1,2*/    
merge_router #(
    .input_mask                     (input_mask_1_2),
    .output_sel                     (output_sel_1_2)
)router11(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_1_2),
    .valid_i                        (valid_i_1_2),
    .ready_o                        (ready_o_1_2),
    .data_o                         (data_o_1_2),
    .valid_o                        (valid_o_1_2),
    .ready_i                        (ready_i_1_2)
);


always@(*) begin
    data_i_1_2[3] = data_o_1_1[4];
    valid_i_1_2[3] = valid_o_1_1[4];
    ready_i_1_2[3] = ready_o_1_1[4];
    data_i_1_2[4] = data_o_1_3[3];
    valid_i_1_2[4] = valid_o_1_3[3];
    ready_i_1_2[4] = ready_o_1_3[3];
    data_i_1_2[1] = data_o_0_2[2];
    valid_i_1_2[1] = valid_o_0_2[2];
    ready_i_1_2[1] = ready_o_0_2[2];
    data_i_1_2[2] = data_o_2_2[1];
    valid_i_1_2[2] = valid_o_2_2[1];
    ready_i_1_2[2] = ready_o_2_2[1];
    data_i_1_2[0] = data_i[1][2];
    valid_i_1_2[0] = valid_i[1][2];
    ready_i_1_2[0] = ready_i[1][2];
end


/*Router 1,3*/    
merge_router #(
    .input_mask                     (input_mask_1_3),
    .output_sel                     (output_sel_1_3)
)router16(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_1_3),
    .valid_i                        (valid_i_1_3),
    .ready_o                        (ready_o_1_3),
    .data_o                         (data_o_1_3),
    .valid_o                        (valid_o_1_3),
    .ready_i                        (ready_i_1_3)
);


always@(*) begin
    data_i_1_3[3] = data_o_1_2[4];
    valid_i_1_3[3] = valid_o_1_2[4];
    ready_i_1_3[3] = ready_o_1_2[4];
    data_i_1_3[4] = data_o_1_4[3];
    valid_i_1_3[4] = valid_o_1_4[3];
    ready_i_1_3[4] = ready_o_1_4[3];
    data_i_1_3[1] = data_o_0_3[2];
    valid_i_1_3[1] = valid_o_0_3[2];
    ready_i_1_3[1] = ready_o_0_3[2];
    data_i_1_3[2] = data_o_2_3[1];
    valid_i_1_3[2] = valid_o_2_3[1];
    ready_i_1_3[2] = ready_o_2_3[1];
    data_i_1_3[0] = data_i[1][3];
    valid_i_1_3[0] = valid_i[1][3];
    ready_i_1_3[0] = ready_i[1][3];
end


/*Router 1,4*/    
merge_router #(
    .input_mask                     (input_mask_1_4),
    .output_sel                     (output_sel_1_4)
)router21(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_1_4),
    .valid_i                        (valid_i_1_4),
    .ready_o                        (ready_o_1_4),
    .data_o                         (data_o_1_4),
    .valid_o                        (valid_o_1_4),
    .ready_i                        (ready_i_1_4)
);


always@(*) begin
    data_i_1_4[3] = data_o_1_3[4];
    valid_i_1_4[3] = valid_o_1_3[4];
    ready_i_1_4[3] = ready_o_1_3[4];
    data_i_1_4[4] = data_o_1_5[3];
    valid_i_1_4[4] = valid_o_1_5[3];
    ready_i_1_4[4] = ready_o_1_5[3];
    data_i_1_4[1] = data_o_0_4[2];
    valid_i_1_4[1] = valid_o_0_4[2];
    ready_i_1_4[1] = ready_o_0_4[2];
    data_i_1_4[2] = data_o_2_4[1];
    valid_i_1_4[2] = valid_o_2_4[1];
    ready_i_1_4[2] = ready_o_2_4[1];
    data_i_1_4[0] = data_i[1][4];
    valid_i_1_4[0] = valid_i[1][4];
    ready_i_1_4[0] = ready_i[1][4];
end


/*Router 1,5*/    
merge_router #(
    .input_mask                     (input_mask_1_5),
    .output_sel                     (output_sel_1_5)
)router26(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_1_5),
    .valid_i                        (valid_i_1_5),
    .ready_o                        (ready_o_1_5),
    .data_o                         (data_o_1_5),
    .valid_o                        (valid_o_1_5),
    .ready_i                        (ready_i_1_5)
);


always@(*) begin
    data_i_1_5[3] = data_o_1_4[4];
    valid_i_1_5[3] = valid_o_1_4[4];
    ready_i_1_5[3] = ready_o_1_4[4];
    data_i_1_5[1] = data_o_0_5[2];
    valid_i_1_5[1] = valid_o_0_5[2];
    ready_i_1_5[1] = ready_o_0_5[2];
    data_i_1_5[2] = data_o_2_5[1];
    valid_i_1_5[2] = valid_o_2_5[1];
    ready_i_1_5[2] = ready_o_2_5[1];
    data_i_1_5[0] = data_i[1][5];
    valid_i_1_5[0] = valid_i[1][5];
    ready_i_1_5[0] = ready_i[1][5];
end


/*Router 2,0*/    
merge_router #(
    .input_mask                     (input_mask_2_0),
    .output_sel                     (output_sel_2_0)
)router2(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_2_0),
    .valid_i                        (valid_i_2_0),
    .ready_o                        (ready_o_2_0),
    .data_o                         (data_o_2_0),
    .valid_o                        (valid_o_2_0),
    .ready_i                        (ready_i_2_0)
);


always@(*) begin
    data_i_2_0[4] = data_o_2_1[3];
    valid_i_2_0[4] = valid_o_2_1[3];
    ready_i_2_0[4] = ready_o_2_1[3];
    data_i_2_0[1] = data_o_1_0[2];
    valid_i_2_0[1] = valid_o_1_0[2];
    ready_i_2_0[1] = ready_o_1_0[2];
    data_i_2_0[2] = data_o_3_0[1];
    valid_i_2_0[2] = valid_o_3_0[1];
    ready_i_2_0[2] = ready_o_3_0[1];
    data_i_2_0[0] = data_i[2][0];
    valid_i_2_0[0] = valid_i[2][0];
    ready_i_2_0[0] = ready_i[2][0];
end


/*Router 2,1*/    
merge_router #(
    .input_mask                     (input_mask_2_1),
    .output_sel                     (output_sel_2_1)
)router7(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_2_1),
    .valid_i                        (valid_i_2_1),
    .ready_o                        (ready_o_2_1),
    .data_o                         (data_o_2_1),
    .valid_o                        (valid_o_2_1),
    .ready_i                        (ready_i_2_1)
);


always@(*) begin
    data_i_2_1[3] = data_o_2_0[4];
    valid_i_2_1[3] = valid_o_2_0[4];
    ready_i_2_1[3] = ready_o_2_0[4];
    data_i_2_1[4] = data_o_2_2[3];
    valid_i_2_1[4] = valid_o_2_2[3];
    ready_i_2_1[4] = ready_o_2_2[3];
    data_i_2_1[1] = data_o_1_1[2];
    valid_i_2_1[1] = valid_o_1_1[2];
    ready_i_2_1[1] = ready_o_1_1[2];
    data_i_2_1[2] = data_o_3_1[1];
    valid_i_2_1[2] = valid_o_3_1[1];
    ready_i_2_1[2] = ready_o_3_1[1];
    data_i_2_1[0] = data_i[2][1];
    valid_i_2_1[0] = valid_i[2][1];
    ready_i_2_1[0] = ready_i[2][1];
end


/*Router 2,2*/    
merge_router #(
    .input_mask                     (input_mask_2_2),
    .output_sel                     (output_sel_2_2)
)router12(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_2_2),
    .valid_i                        (valid_i_2_2),
    .ready_o                        (ready_o_2_2),
    .data_o                         (data_o_2_2),
    .valid_o                        (valid_o_2_2),
    .ready_i                        (ready_i_2_2)
);


always@(*) begin
    data_i_2_2[3] = data_o_2_1[4];
    valid_i_2_2[3] = valid_o_2_1[4];
    ready_i_2_2[3] = ready_o_2_1[4];
    data_i_2_2[4] = data_o_2_3[3];
    valid_i_2_2[4] = valid_o_2_3[3];
    ready_i_2_2[4] = ready_o_2_3[3];
    data_i_2_2[1] = data_o_1_2[2];
    valid_i_2_2[1] = valid_o_1_2[2];
    ready_i_2_2[1] = ready_o_1_2[2];
    data_i_2_2[2] = data_o_3_2[1];
    valid_i_2_2[2] = valid_o_3_2[1];
    ready_i_2_2[2] = ready_o_3_2[1];
    data_i_2_2[0] = data_i[2][2];
    valid_i_2_2[0] = valid_i[2][2];
    ready_i_2_2[0] = ready_i[2][2];
end


/*Router 2,3*/    
merge_router #(
    .input_mask                     (input_mask_2_3),
    .output_sel                     (output_sel_2_3)
)router17(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_2_3),
    .valid_i                        (valid_i_2_3),
    .ready_o                        (ready_o_2_3),
    .data_o                         (data_o_2_3),
    .valid_o                        (valid_o_2_3),
    .ready_i                        (ready_i_2_3)
);


always@(*) begin
    data_i_2_3[3] = data_o_2_2[4];
    valid_i_2_3[3] = valid_o_2_2[4];
    ready_i_2_3[3] = ready_o_2_2[4];
    data_i_2_3[4] = data_o_2_4[3];
    valid_i_2_3[4] = valid_o_2_4[3];
    ready_i_2_3[4] = ready_o_2_4[3];
    data_i_2_3[1] = data_o_1_3[2];
    valid_i_2_3[1] = valid_o_1_3[2];
    ready_i_2_3[1] = ready_o_1_3[2];
    data_i_2_3[2] = data_o_3_3[1];
    valid_i_2_3[2] = valid_o_3_3[1];
    ready_i_2_3[2] = ready_o_3_3[1];
    data_i_2_3[0] = data_i[2][3];
    valid_i_2_3[0] = valid_i[2][3];
    ready_i_2_3[0] = ready_i[2][3];
end


/*Router 2,4*/    
merge_router #(
    .input_mask                     (input_mask_2_4),
    .output_sel                     (output_sel_2_4)
)router22(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_2_4),
    .valid_i                        (valid_i_2_4),
    .ready_o                        (ready_o_2_4),
    .data_o                         (data_o_2_4),
    .valid_o                        (valid_o_2_4),
    .ready_i                        (ready_i_2_4)
);


always@(*) begin
    data_i_2_4[3] = data_o_2_3[4];
    valid_i_2_4[3] = valid_o_2_3[4];
    ready_i_2_4[3] = ready_o_2_3[4];
    data_i_2_4[4] = data_o_2_5[3];
    valid_i_2_4[4] = valid_o_2_5[3];
    ready_i_2_4[4] = ready_o_2_5[3];
    data_i_2_4[1] = data_o_1_4[2];
    valid_i_2_4[1] = valid_o_1_4[2];
    ready_i_2_4[1] = ready_o_1_4[2];
    data_i_2_4[2] = data_o_3_4[1];
    valid_i_2_4[2] = valid_o_3_4[1];
    ready_i_2_4[2] = ready_o_3_4[1];
    data_i_2_4[0] = data_i[2][4];
    valid_i_2_4[0] = valid_i[2][4];
    ready_i_2_4[0] = ready_i[2][4];
end


/*Router 2,5*/    
merge_router #(
    .input_mask                     (input_mask_2_5),
    .output_sel                     (output_sel_2_5)
)router27(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_2_5),
    .valid_i                        (valid_i_2_5),
    .ready_o                        (ready_o_2_5),
    .data_o                         (data_o_2_5),
    .valid_o                        (valid_o_2_5),
    .ready_i                        (ready_i_2_5)
);


always@(*) begin
    data_i_2_5[3] = data_o_2_4[4];
    valid_i_2_5[3] = valid_o_2_4[4];
    ready_i_2_5[3] = ready_o_2_4[4];
    data_i_2_5[1] = data_o_1_5[2];
    valid_i_2_5[1] = valid_o_1_5[2];
    ready_i_2_5[1] = ready_o_1_5[2];
    data_i_2_5[2] = data_o_3_5[1];
    valid_i_2_5[2] = valid_o_3_5[1];
    ready_i_2_5[2] = ready_o_3_5[1];
    data_i_2_5[0] = data_i[2][5];
    valid_i_2_5[0] = valid_i[2][5];
    ready_i_2_5[0] = ready_i[2][5];
end


/*Router 3,0*/    
merge_router #(
    .input_mask                     (input_mask_3_0),
    .output_sel                     (output_sel_3_0)
)router3(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_3_0),
    .valid_i                        (valid_i_3_0),
    .ready_o                        (ready_o_3_0),
    .data_o                         (data_o_3_0),
    .valid_o                        (valid_o_3_0),
    .ready_i                        (ready_i_3_0)
);


always@(*) begin
    data_i_3_0[4] = data_o_3_1[3];
    valid_i_3_0[4] = valid_o_3_1[3];
    ready_i_3_0[4] = ready_o_3_1[3];
    data_i_3_0[1] = data_o_2_0[2];
    valid_i_3_0[1] = valid_o_2_0[2];
    ready_i_3_0[1] = ready_o_2_0[2];
    data_i_3_0[2] = data_o_4_0[1];
    valid_i_3_0[2] = valid_o_4_0[1];
    ready_i_3_0[2] = ready_o_4_0[1];
    data_i_3_0[0] = data_i[3][0];
    valid_i_3_0[0] = valid_i[3][0];
    ready_i_3_0[0] = ready_i[3][0];
end


/*Router 3,1*/    
merge_router #(
    .input_mask                     (input_mask_3_1),
    .output_sel                     (output_sel_3_1)
)router8(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_3_1),
    .valid_i                        (valid_i_3_1),
    .ready_o                        (ready_o_3_1),
    .data_o                         (data_o_3_1),
    .valid_o                        (valid_o_3_1),
    .ready_i                        (ready_i_3_1)
);


always@(*) begin
    data_i_3_1[3] = data_o_3_0[4];
    valid_i_3_1[3] = valid_o_3_0[4];
    ready_i_3_1[3] = ready_o_3_0[4];
    data_i_3_1[4] = data_o_3_2[3];
    valid_i_3_1[4] = valid_o_3_2[3];
    ready_i_3_1[4] = ready_o_3_2[3];
    data_i_3_1[1] = data_o_2_1[2];
    valid_i_3_1[1] = valid_o_2_1[2];
    ready_i_3_1[1] = ready_o_2_1[2];
    data_i_3_1[2] = data_o_4_1[1];
    valid_i_3_1[2] = valid_o_4_1[1];
    ready_i_3_1[2] = ready_o_4_1[1];
    data_i_3_1[0] = data_i[3][1];
    valid_i_3_1[0] = valid_i[3][1];
    ready_i_3_1[0] = ready_i[3][1];
end


/*Router 3,2*/    
merge_router #(
    .input_mask                     (input_mask_3_2),
    .output_sel                     (output_sel_3_2)
)router13(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_3_2),
    .valid_i                        (valid_i_3_2),
    .ready_o                        (ready_o_3_2),
    .data_o                         (data_o_3_2),
    .valid_o                        (valid_o_3_2),
    .ready_i                        (ready_i_3_2)
);


always@(*) begin
    data_i_3_2[3] = data_o_3_1[4];
    valid_i_3_2[3] = valid_o_3_1[4];
    ready_i_3_2[3] = ready_o_3_1[4];
    data_i_3_2[4] = data_o_3_3[3];
    valid_i_3_2[4] = valid_o_3_3[3];
    ready_i_3_2[4] = ready_o_3_3[3];
    data_i_3_2[1] = data_o_2_2[2];
    valid_i_3_2[1] = valid_o_2_2[2];
    ready_i_3_2[1] = ready_o_2_2[2];
    data_i_3_2[2] = data_o_4_2[1];
    valid_i_3_2[2] = valid_o_4_2[1];
    ready_i_3_2[2] = ready_o_4_2[1];
    data_i_3_2[0] = data_i[3][2];
    valid_i_3_2[0] = valid_i[3][2];
    ready_i_3_2[0] = ready_i[3][2];
end


/*Router 3,3*/    
merge_router #(
    .input_mask                     (input_mask_3_3),
    .output_sel                     (output_sel_3_3)
)router18(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_3_3),
    .valid_i                        (valid_i_3_3),
    .ready_o                        (ready_o_3_3),
    .data_o                         (data_o_3_3),
    .valid_o                        (valid_o_3_3),
    .ready_i                        (ready_i_3_3)
);


always@(*) begin
    data_i_3_3[3] = data_o_3_2[4];
    valid_i_3_3[3] = valid_o_3_2[4];
    ready_i_3_3[3] = ready_o_3_2[4];
    data_i_3_3[4] = data_o_3_4[3];
    valid_i_3_3[4] = valid_o_3_4[3];
    ready_i_3_3[4] = ready_o_3_4[3];
    data_i_3_3[1] = data_o_2_3[2];
    valid_i_3_3[1] = valid_o_2_3[2];
    ready_i_3_3[1] = ready_o_2_3[2];
    data_i_3_3[2] = data_o_4_3[1];
    valid_i_3_3[2] = valid_o_4_3[1];
    ready_i_3_3[2] = ready_o_4_3[1];
    data_i_3_3[0] = data_i[3][3];
    valid_i_3_3[0] = valid_i[3][3];
    ready_i_3_3[0] = ready_i[3][3];
end


/*Router 3,4*/    
merge_router #(
    .input_mask                     (input_mask_3_4),
    .output_sel                     (output_sel_3_4)
)router23(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_3_4),
    .valid_i                        (valid_i_3_4),
    .ready_o                        (ready_o_3_4),
    .data_o                         (data_o_3_4),
    .valid_o                        (valid_o_3_4),
    .ready_i                        (ready_i_3_4)
);


always@(*) begin
    data_i_3_4[3] = data_o_3_3[4];
    valid_i_3_4[3] = valid_o_3_3[4];
    ready_i_3_4[3] = ready_o_3_3[4];
    data_i_3_4[4] = data_o_3_5[3];
    valid_i_3_4[4] = valid_o_3_5[3];
    ready_i_3_4[4] = ready_o_3_5[3];
    data_i_3_4[1] = data_o_2_4[2];
    valid_i_3_4[1] = valid_o_2_4[2];
    ready_i_3_4[1] = ready_o_2_4[2];
    data_i_3_4[2] = data_o_4_4[1];
    valid_i_3_4[2] = valid_o_4_4[1];
    ready_i_3_4[2] = ready_o_4_4[1];
    data_i_3_4[0] = data_i[3][4];
    valid_i_3_4[0] = valid_i[3][4];
    ready_i_3_4[0] = ready_i[3][4];
end


/*Router 3,5*/    
merge_router #(
    .input_mask                     (input_mask_3_5),
    .output_sel                     (output_sel_3_5)
)router28(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_3_5),
    .valid_i                        (valid_i_3_5),
    .ready_o                        (ready_o_3_5),
    .data_o                         (data_o_3_5),
    .valid_o                        (valid_o_3_5),
    .ready_i                        (ready_i_3_5)
);


always@(*) begin
    data_i_3_5[3] = data_o_3_4[4];
    valid_i_3_5[3] = valid_o_3_4[4];
    ready_i_3_5[3] = ready_o_3_4[4];
    data_i_3_5[1] = data_o_2_5[2];
    valid_i_3_5[1] = valid_o_2_5[2];
    ready_i_3_5[1] = ready_o_2_5[2];
    data_i_3_5[2] = data_o_4_5[1];
    valid_i_3_5[2] = valid_o_4_5[1];
    ready_i_3_5[2] = ready_o_4_5[1];
    data_i_3_5[0] = data_i[3][5];
    valid_i_3_5[0] = valid_i[3][5];
    ready_i_3_5[0] = ready_i[3][5];
end


/*Router 4,0*/    
merge_router #(
    .input_mask                     (input_mask_4_0),
    .output_sel                     (output_sel_4_0)
)router4(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_4_0),
    .valid_i                        (valid_i_4_0),
    .ready_o                        (ready_o_4_0),
    .data_o                         (data_o_4_0),
    .valid_o                        (valid_o_4_0),
    .ready_i                        (ready_i_4_0)
);


always@(*) begin
    data_i_4_0[4] = data_o_4_1[3];
    valid_i_4_0[4] = valid_o_4_1[3];
    ready_i_4_0[4] = ready_o_4_1[3];
    data_i_4_0[1] = data_o_3_0[2];
    valid_i_4_0[1] = valid_o_3_0[2];
    ready_i_4_0[1] = ready_o_3_0[2];
    data_i_4_0[0] = data_i[4][0];
    valid_i_4_0[0] = valid_i[4][0];
    ready_i_4_0[0] = ready_i[4][0];
end


/*Router 4,1*/    
merge_router #(
    .input_mask                     (input_mask_4_1),
    .output_sel                     (output_sel_4_1)
)router9(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_4_1),
    .valid_i                        (valid_i_4_1),
    .ready_o                        (ready_o_4_1),
    .data_o                         (data_o_4_1),
    .valid_o                        (valid_o_4_1),
    .ready_i                        (ready_i_4_1)
);


always@(*) begin
    data_i_4_1[3] = data_o_4_0[4];
    valid_i_4_1[3] = valid_o_4_0[4];
    ready_i_4_1[3] = ready_o_4_0[4];
    data_i_4_1[4] = data_o_4_2[3];
    valid_i_4_1[4] = valid_o_4_2[3];
    ready_i_4_1[4] = ready_o_4_2[3];
    data_i_4_1[1] = data_o_3_1[2];
    valid_i_4_1[1] = valid_o_3_1[2];
    ready_i_4_1[1] = ready_o_3_1[2];
    data_i_4_1[0] = data_i[4][1];
    valid_i_4_1[0] = valid_i[4][1];
    ready_i_4_1[0] = ready_i[4][1];
end


/*Router 4,2*/    
merge_router #(
    .input_mask                     (input_mask_4_2),
    .output_sel                     (output_sel_4_2)
)router14(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_4_2),
    .valid_i                        (valid_i_4_2),
    .ready_o                        (ready_o_4_2),
    .data_o                         (data_o_4_2),
    .valid_o                        (valid_o_4_2),
    .ready_i                        (ready_i_4_2)
);


always@(*) begin
    data_i_4_2[3] = data_o_4_1[4];
    valid_i_4_2[3] = valid_o_4_1[4];
    ready_i_4_2[3] = ready_o_4_1[4];
    data_i_4_2[4] = data_o_4_3[3];
    valid_i_4_2[4] = valid_o_4_3[3];
    ready_i_4_2[4] = ready_o_4_3[3];
    data_i_4_2[1] = data_o_3_2[2];
    valid_i_4_2[1] = valid_o_3_2[2];
    ready_i_4_2[1] = ready_o_3_2[2];
    data_i_4_2[0] = data_i[4][2];
    valid_i_4_2[0] = valid_i[4][2];
    ready_i_4_2[0] = ready_i[4][2];
end


/*Router 4,3*/    
merge_router #(
    .input_mask                     (input_mask_4_3),
    .output_sel                     (output_sel_4_3)
)router19(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_4_3),
    .valid_i                        (valid_i_4_3),
    .ready_o                        (ready_o_4_3),
    .data_o                         (data_o_4_3),
    .valid_o                        (valid_o_4_3),
    .ready_i                        (ready_i_4_3)
);


always@(*) begin
    data_i_4_3[3] = data_o_4_2[4];
    valid_i_4_3[3] = valid_o_4_2[4];
    ready_i_4_3[3] = ready_o_4_2[4];
    data_i_4_3[4] = data_o_4_4[3];
    valid_i_4_3[4] = valid_o_4_4[3];
    ready_i_4_3[4] = ready_o_4_4[3];
    data_i_4_3[1] = data_o_3_3[2];
    valid_i_4_3[1] = valid_o_3_3[2];
    ready_i_4_3[1] = ready_o_3_3[2];
    data_i_4_3[0] = data_i[4][3];
    valid_i_4_3[0] = valid_i[4][3];
    ready_i_4_3[0] = ready_i[4][3];
end


/*Router 4,4*/    
merge_router #(
    .input_mask                     (input_mask_4_4),
    .output_sel                     (output_sel_4_4)
)router24(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_4_4),
    .valid_i                        (valid_i_4_4),
    .ready_o                        (ready_o_4_4),
    .data_o                         (data_o_4_4),
    .valid_o                        (valid_o_4_4),
    .ready_i                        (ready_i_4_4)
);


always@(*) begin
    data_i_4_4[3] = data_o_4_3[4];
    valid_i_4_4[3] = valid_o_4_3[4];
    ready_i_4_4[3] = ready_o_4_3[4];
    data_i_4_4[4] = data_o_4_5[3];
    valid_i_4_4[4] = valid_o_4_5[3];
    ready_i_4_4[4] = ready_o_4_5[3];
    data_i_4_4[1] = data_o_3_4[2];
    valid_i_4_4[1] = valid_o_3_4[2];
    ready_i_4_4[1] = ready_o_3_4[2];
    data_i_4_4[0] = data_i[4][4];
    valid_i_4_4[0] = valid_i[4][4];
    ready_i_4_4[0] = ready_i[4][4];
end


/*Router 4,5*/    
merge_router #(
    .input_mask                     (input_mask_4_5),
    .output_sel                     (output_sel_4_5)
)router29(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_4_5),
    .valid_i                        (valid_i_4_5),
    .ready_o                        (ready_o_4_5),
    .data_o                         (data_o_4_5),
    .valid_o                        (valid_o_4_5),
    .ready_i                        (ready_i_4_5)
);


always@(*) begin
    data_i_4_5[3] = data_o_4_4[4];
    valid_i_4_5[3] = valid_o_4_4[4];
    ready_i_4_5[3] = ready_o_4_4[4];
    data_i_4_5[1] = data_o_3_5[2];
    valid_i_4_5[1] = valid_o_3_5[2];
    ready_i_4_5[1] = ready_o_3_5[2];
    data_i_4_5[0] = data_i[4][5];
    valid_i_4_5[0] = valid_i[4][5];
    ready_i_4_5[0] = ready_i[4][5];
end


endmodule
