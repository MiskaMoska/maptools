
`ifndef __MERGE_NETWORK_CONFIG_SVH_
`define __MERGE_NETWORK_CONFIG_SVH_
    
localparam input_mask_0_0 = 5'b10000;
localparam output_sel_0_0 = 5'b00000;
localparam input_mask_0_1 = 5'b10000;
localparam output_sel_0_1 = 5'b00000;
localparam input_mask_0_2 = 5'b10000;
localparam output_sel_0_2 = 5'b00000;
localparam input_mask_0_3 = 5'b00100;
localparam output_sel_0_3 = 5'b10000;
localparam input_mask_0_4 = 5'b10000;
localparam output_sel_0_4 = 5'b00100;
localparam input_mask_0_5 = 5'b10000;
localparam output_sel_0_5 = 5'b00100;
localparam input_mask_0_6 = 5'b10000;
localparam output_sel_0_6 = 5'b00100;
localparam input_mask_0_7 = 5'b10000;
localparam output_sel_0_7 = 5'b00001;
localparam input_mask_0_8 = 5'b10010;
localparam output_sel_0_8 = 5'b00100;
localparam input_mask_0_9 = 5'b10000;
localparam output_sel_0_9 = 5'b00100;
localparam input_mask_0_10 = 5'b10000;
localparam output_sel_0_10 = 5'b00100;
localparam input_mask_0_11 = 5'b10000;
localparam output_sel_0_11 = 5'b00100;
localparam input_mask_0_12 = 5'b10000;
localparam output_sel_0_12 = 5'b00100;
localparam input_mask_0_13 = 5'b10000;
localparam output_sel_0_13 = 5'b00100;
localparam input_mask_0_14 = 5'b10000;
localparam output_sel_0_14 = 5'b00100;
localparam input_mask_0_15 = 5'b10000;
localparam output_sel_0_15 = 5'b00100;
localparam input_mask_0_16 = 5'b10000;
localparam output_sel_0_16 = 5'b00100;
localparam input_mask_0_17 = 5'b10000;
localparam output_sel_0_17 = 5'b00001;
localparam input_mask_0_18 = 5'b10010;
localparam output_sel_0_18 = 5'b00100;
localparam input_mask_0_19 = 5'b10000;
localparam output_sel_0_19 = 5'b00100;
localparam input_mask_0_20 = 5'b10000;
localparam output_sel_0_20 = 5'b00100;
localparam input_mask_0_21 = 5'b10000;
localparam output_sel_0_21 = 5'b00100;
localparam input_mask_0_22 = 5'b10000;
localparam output_sel_0_22 = 5'b00100;
localparam input_mask_0_23 = 5'b00100;
localparam output_sel_0_23 = 5'b10000;
localparam input_mask_0_24 = 5'b10000;
localparam output_sel_0_24 = 5'b00100;
localparam input_mask_1_0 = 5'b10000;
localparam output_sel_1_0 = 5'b00000;
localparam input_mask_1_1 = 5'b10000;
localparam output_sel_1_1 = 5'b00100;
localparam input_mask_1_2 = 5'b10000;
localparam output_sel_1_2 = 5'b00000;
localparam input_mask_1_3 = 5'b10000;
localparam output_sel_1_3 = 5'b01000;
localparam input_mask_1_4 = 5'b01000;
localparam output_sel_1_4 = 5'b10000;
localparam input_mask_1_5 = 5'b11000;
localparam output_sel_1_5 = 5'b00001;
localparam input_mask_1_6 = 5'b01010;
localparam output_sel_1_6 = 5'b10000;
localparam input_mask_1_7 = 5'b10000;
localparam output_sel_1_7 = 5'b00001;
localparam input_mask_1_8 = 5'b01010;
localparam output_sel_1_8 = 5'b10000;
localparam input_mask_1_9 = 5'b11000;
localparam output_sel_1_9 = 5'b00001;
localparam input_mask_1_10 = 5'b01010;
localparam output_sel_1_10 = 5'b10000;
localparam input_mask_1_11 = 5'b11000;
localparam output_sel_1_11 = 5'b00001;
localparam input_mask_1_12 = 5'b01010;
localparam output_sel_1_12 = 5'b10000;
localparam input_mask_1_13 = 5'b11000;
localparam output_sel_1_13 = 5'b00001;
localparam input_mask_1_14 = 5'b01010;
localparam output_sel_1_14 = 5'b10000;
localparam input_mask_1_15 = 5'b01000;
localparam output_sel_1_15 = 5'b10000;
localparam input_mask_1_16 = 5'b01000;
localparam output_sel_1_16 = 5'b10000;
localparam input_mask_1_17 = 5'b10000;
localparam output_sel_1_17 = 5'b00001;
localparam input_mask_1_18 = 5'b01010;
localparam output_sel_1_18 = 5'b10000;
localparam input_mask_1_19 = 5'b01000;
localparam output_sel_1_19 = 5'b10000;
localparam input_mask_1_20 = 5'b01000;
localparam output_sel_1_20 = 5'b10000;
localparam input_mask_1_21 = 5'b11000;
localparam output_sel_1_21 = 5'b00001;
localparam input_mask_1_22 = 5'b01010;
localparam output_sel_1_22 = 5'b10000;
localparam input_mask_1_23 = 5'b10000;
localparam output_sel_1_23 = 5'b01000;
localparam input_mask_1_24 = 5'b01000;
localparam output_sel_1_24 = 5'b10000;
localparam input_mask_2_0 = 5'b10000;
localparam output_sel_2_0 = 5'b00000;
localparam input_mask_2_1 = 5'b01000;
localparam output_sel_2_1 = 5'b10000;
localparam input_mask_2_2 = 5'b10000;
localparam output_sel_2_2 = 5'b00100;
localparam input_mask_2_3 = 5'b00100;
localparam output_sel_2_3 = 5'b10000;
localparam input_mask_2_4 = 5'b10000;
localparam output_sel_2_4 = 5'b00100;
localparam input_mask_2_5 = 5'b10000;
localparam output_sel_2_5 = 5'b00000;
localparam input_mask_2_6 = 5'b10000;
localparam output_sel_2_6 = 5'b00100;
localparam input_mask_2_7 = 5'b10000;
localparam output_sel_2_7 = 5'b00000;
localparam input_mask_2_8 = 5'b10000;
localparam output_sel_2_8 = 5'b00100;
localparam input_mask_2_9 = 5'b10000;
localparam output_sel_2_9 = 5'b00000;
localparam input_mask_2_10 = 5'b10000;
localparam output_sel_2_10 = 5'b00100;
localparam input_mask_2_11 = 5'b00100;
localparam output_sel_2_11 = 5'b10000;
localparam input_mask_2_12 = 5'b10000;
localparam output_sel_2_12 = 5'b00100;
localparam input_mask_2_13 = 5'b10000;
localparam output_sel_2_13 = 5'b00100;
localparam input_mask_2_14 = 5'b10000;
localparam output_sel_2_14 = 5'b00100;
localparam input_mask_2_15 = 5'b10000;
localparam output_sel_2_15 = 5'b00100;
localparam input_mask_2_16 = 5'b10000;
localparam output_sel_2_16 = 5'b00100;
localparam input_mask_2_17 = 5'b10000;
localparam output_sel_2_17 = 5'b00100;
localparam input_mask_2_18 = 5'b10000;
localparam output_sel_2_18 = 5'b00100;
localparam input_mask_2_19 = 5'b10000;
localparam output_sel_2_19 = 5'b00100;
localparam input_mask_2_20 = 5'b10000;
localparam output_sel_2_20 = 5'b00100;
localparam input_mask_2_21 = 5'b10000;
localparam output_sel_2_21 = 5'b00100;
localparam input_mask_2_22 = 5'b10000;
localparam output_sel_2_22 = 5'b00100;
localparam input_mask_2_23 = 5'b10000;
localparam output_sel_2_23 = 5'b00100;
localparam input_mask_2_24 = 5'b10000;
localparam output_sel_2_24 = 5'b00000;
localparam input_mask_3_0 = 5'b10000;
localparam output_sel_3_0 = 5'b00000;
localparam input_mask_3_1 = 5'b10000;
localparam output_sel_3_1 = 5'b00000;
localparam input_mask_3_2 = 5'b01000;
localparam output_sel_3_2 = 5'b10000;
localparam input_mask_3_3 = 5'b10000;
localparam output_sel_3_3 = 5'b01000;
localparam input_mask_3_4 = 5'b01000;
localparam output_sel_3_4 = 5'b10000;
localparam input_mask_3_5 = 5'b10000;
localparam output_sel_3_5 = 5'b00000;
localparam input_mask_3_6 = 5'b01000;
localparam output_sel_3_6 = 5'b10000;
localparam input_mask_3_7 = 5'b10000;
localparam output_sel_3_7 = 5'b00000;
localparam input_mask_3_8 = 5'b01000;
localparam output_sel_3_8 = 5'b10000;
localparam input_mask_3_9 = 5'b10000;
localparam output_sel_3_9 = 5'b00000;
localparam input_mask_3_10 = 5'b11000;
localparam output_sel_3_10 = 5'b00100;
localparam input_mask_3_11 = 5'b10100;
localparam output_sel_3_11 = 5'b01000;
localparam input_mask_3_12 = 5'b11000;
localparam output_sel_3_12 = 5'b00100;
localparam input_mask_3_13 = 5'b01100;
localparam output_sel_3_13 = 5'b10000;
localparam input_mask_3_14 = 5'b11000;
localparam output_sel_3_14 = 5'b00100;
localparam input_mask_3_15 = 5'b01000;
localparam output_sel_3_15 = 5'b10000;
localparam input_mask_3_16 = 5'b11000;
localparam output_sel_3_16 = 5'b00100;
localparam input_mask_3_17 = 5'b11000;
localparam output_sel_3_17 = 5'b00100;
localparam input_mask_3_18 = 5'b11000;
localparam output_sel_3_18 = 5'b00100;
localparam input_mask_3_19 = 5'b01000;
localparam output_sel_3_19 = 5'b10000;
localparam input_mask_3_20 = 5'b11000;
localparam output_sel_3_20 = 5'b00100;
localparam input_mask_3_21 = 5'b11000;
localparam output_sel_3_21 = 5'b00100;
localparam input_mask_3_22 = 5'b11000;
localparam output_sel_3_22 = 5'b00100;
localparam input_mask_3_23 = 5'b01000;
localparam output_sel_3_23 = 5'b10000;
localparam input_mask_3_24 = 5'b10000;
localparam output_sel_3_24 = 5'b00000;
localparam input_mask_4_0 = 5'b10000;
localparam output_sel_4_0 = 5'b00000;
localparam input_mask_4_1 = 5'b10000;
localparam output_sel_4_1 = 5'b00000;
localparam input_mask_4_2 = 5'b10000;
localparam output_sel_4_2 = 5'b00000;
localparam input_mask_4_3 = 5'b00100;
localparam output_sel_4_3 = 5'b10000;
localparam input_mask_4_4 = 5'b10000;
localparam output_sel_4_4 = 5'b00000;
localparam input_mask_4_5 = 5'b10000;
localparam output_sel_4_5 = 5'b00000;
localparam input_mask_4_6 = 5'b10000;
localparam output_sel_4_6 = 5'b00000;
localparam input_mask_4_7 = 5'b10000;
localparam output_sel_4_7 = 5'b00000;
localparam input_mask_4_8 = 5'b10000;
localparam output_sel_4_8 = 5'b00000;
localparam input_mask_4_9 = 5'b10000;
localparam output_sel_4_9 = 5'b00000;
localparam input_mask_4_10 = 5'b11000;
localparam output_sel_4_10 = 5'b00100;
localparam input_mask_4_11 = 5'b10100;
localparam output_sel_4_11 = 5'b01000;
localparam input_mask_4_12 = 5'b11000;
localparam output_sel_4_12 = 5'b00100;
localparam input_mask_4_13 = 5'b10100;
localparam output_sel_4_13 = 5'b01000;
localparam input_mask_4_14 = 5'b11000;
localparam output_sel_4_14 = 5'b00100;
localparam input_mask_4_15 = 5'b00100;
localparam output_sel_4_15 = 5'b10000;
localparam input_mask_4_16 = 5'b11000;
localparam output_sel_4_16 = 5'b00100;
localparam input_mask_4_17 = 5'b11000;
localparam output_sel_4_17 = 5'b00100;
localparam input_mask_4_18 = 5'b11000;
localparam output_sel_4_18 = 5'b00100;
localparam input_mask_4_19 = 5'b10000;
localparam output_sel_4_19 = 5'b00100;
localparam input_mask_4_20 = 5'b11000;
localparam output_sel_4_20 = 5'b00100;
localparam input_mask_4_21 = 5'b11000;
localparam output_sel_4_21 = 5'b00100;
localparam input_mask_4_22 = 5'b11000;
localparam output_sel_4_22 = 5'b00100;
localparam input_mask_4_23 = 5'b10000;
localparam output_sel_4_23 = 5'b00100;
localparam input_mask_4_24 = 5'b10000;
localparam output_sel_4_24 = 5'b00000;
localparam input_mask_5_0 = 5'b10000;
localparam output_sel_5_0 = 5'b00000;
localparam input_mask_5_1 = 5'b10000;
localparam output_sel_5_1 = 5'b00000;
localparam input_mask_5_2 = 5'b10000;
localparam output_sel_5_2 = 5'b00000;
localparam input_mask_5_3 = 5'b10000;
localparam output_sel_5_3 = 5'b01000;
localparam input_mask_5_4 = 5'b10000;
localparam output_sel_5_4 = 5'b00000;
localparam input_mask_5_5 = 5'b10000;
localparam output_sel_5_5 = 5'b00000;
localparam input_mask_5_6 = 5'b10000;
localparam output_sel_5_6 = 5'b00000;
localparam input_mask_5_7 = 5'b10000;
localparam output_sel_5_7 = 5'b00000;
localparam input_mask_5_8 = 5'b10000;
localparam output_sel_5_8 = 5'b00000;
localparam input_mask_5_9 = 5'b10000;
localparam output_sel_5_9 = 5'b00000;
localparam input_mask_5_10 = 5'b01000;
localparam output_sel_5_10 = 5'b10000;
localparam input_mask_5_11 = 5'b10000;
localparam output_sel_5_11 = 5'b01000;
localparam input_mask_5_12 = 5'b01000;
localparam output_sel_5_12 = 5'b10000;
localparam input_mask_5_13 = 5'b10000;
localparam output_sel_5_13 = 5'b01000;
localparam input_mask_5_14 = 5'b01000;
localparam output_sel_5_14 = 5'b10000;
localparam input_mask_5_15 = 5'b10000;
localparam output_sel_5_15 = 5'b01000;
localparam input_mask_5_16 = 5'b11000;
localparam output_sel_5_16 = 5'b00100;
localparam input_mask_5_17 = 5'b11000;
localparam output_sel_5_17 = 5'b00100;
localparam input_mask_5_18 = 5'b01000;
localparam output_sel_5_18 = 5'b10000;
localparam input_mask_5_19 = 5'b01000;
localparam output_sel_5_19 = 5'b10000;
localparam input_mask_5_20 = 5'b11000;
localparam output_sel_5_20 = 5'b00100;
localparam input_mask_5_21 = 5'b01100;
localparam output_sel_5_21 = 5'b10000;
localparam input_mask_5_22 = 5'b01000;
localparam output_sel_5_22 = 5'b10000;
localparam input_mask_5_23 = 5'b01000;
localparam output_sel_5_23 = 5'b10000;
localparam input_mask_5_24 = 5'b10000;
localparam output_sel_5_24 = 5'b00000;
localparam input_mask_6_0 = 5'b10000;
localparam output_sel_6_0 = 5'b00000;
localparam input_mask_6_1 = 5'b10000;
localparam output_sel_6_1 = 5'b00000;
localparam input_mask_6_2 = 5'b10000;
localparam output_sel_6_2 = 5'b00000;
localparam input_mask_6_3 = 5'b00100;
localparam output_sel_6_3 = 5'b10000;
localparam input_mask_6_4 = 5'b10000;
localparam output_sel_6_4 = 5'b00000;
localparam input_mask_6_5 = 5'b00100;
localparam output_sel_6_5 = 5'b10000;
localparam input_mask_6_6 = 5'b10000;
localparam output_sel_6_6 = 5'b00000;
localparam input_mask_6_7 = 5'b10000;
localparam output_sel_6_7 = 5'b00100;
localparam input_mask_6_8 = 5'b10000;
localparam output_sel_6_8 = 5'b00000;
localparam input_mask_6_9 = 5'b00100;
localparam output_sel_6_9 = 5'b10000;
localparam input_mask_6_10 = 5'b10000;
localparam output_sel_6_10 = 5'b00100;
localparam input_mask_6_11 = 5'b10000;
localparam output_sel_6_11 = 5'b00100;
localparam input_mask_6_12 = 5'b10000;
localparam output_sel_6_12 = 5'b00100;
localparam input_mask_6_13 = 5'b10000;
localparam output_sel_6_13 = 5'b00100;
localparam input_mask_6_14 = 5'b10000;
localparam output_sel_6_14 = 5'b00100;
localparam input_mask_6_15 = 5'b00100;
localparam output_sel_6_15 = 5'b10000;
localparam input_mask_6_16 = 5'b11000;
localparam output_sel_6_16 = 5'b00100;
localparam input_mask_6_17 = 5'b01100;
localparam output_sel_6_17 = 5'b10000;
localparam input_mask_6_18 = 5'b10000;
localparam output_sel_6_18 = 5'b00100;
localparam input_mask_6_19 = 5'b00100;
localparam output_sel_6_19 = 5'b10000;
localparam input_mask_6_20 = 5'b11000;
localparam output_sel_6_20 = 5'b00100;
localparam input_mask_6_21 = 5'b10100;
localparam output_sel_6_21 = 5'b01000;
localparam input_mask_6_22 = 5'b10000;
localparam output_sel_6_22 = 5'b00100;
localparam input_mask_6_23 = 5'b00100;
localparam output_sel_6_23 = 5'b10000;
localparam input_mask_6_24 = 5'b10000;
localparam output_sel_6_24 = 5'b00000;
localparam input_mask_7_0 = 5'b10000;
localparam output_sel_7_0 = 5'b00000;
localparam input_mask_7_1 = 5'b10000;
localparam output_sel_7_1 = 5'b00000;
localparam input_mask_7_2 = 5'b10000;
localparam output_sel_7_2 = 5'b00100;
localparam input_mask_7_3 = 5'b10000;
localparam output_sel_7_3 = 5'b01000;
localparam input_mask_7_4 = 5'b10000;
localparam output_sel_7_4 = 5'b00000;
localparam input_mask_7_5 = 5'b10000;
localparam output_sel_7_5 = 5'b01000;
localparam input_mask_7_6 = 5'b10000;
localparam output_sel_7_6 = 5'b00000;
localparam input_mask_7_7 = 5'b01000;
localparam output_sel_7_7 = 5'b10000;
localparam input_mask_7_8 = 5'b10000;
localparam output_sel_7_8 = 5'b00000;
localparam input_mask_7_9 = 5'b10000;
localparam output_sel_7_9 = 5'b01000;
localparam input_mask_7_10 = 5'b11000;
localparam output_sel_7_10 = 5'b00100;
localparam input_mask_7_11 = 5'b11000;
localparam output_sel_7_11 = 5'b00100;
localparam input_mask_7_12 = 5'b11000;
localparam output_sel_7_12 = 5'b00100;
localparam input_mask_7_13 = 5'b11000;
localparam output_sel_7_13 = 5'b00100;
localparam input_mask_7_14 = 5'b01000;
localparam output_sel_7_14 = 5'b10000;
localparam input_mask_7_15 = 5'b10000;
localparam output_sel_7_15 = 5'b01000;
localparam input_mask_7_16 = 5'b11000;
localparam output_sel_7_16 = 5'b00100;
localparam input_mask_7_17 = 5'b10100;
localparam output_sel_7_17 = 5'b01000;
localparam input_mask_7_18 = 5'b01000;
localparam output_sel_7_18 = 5'b10000;
localparam input_mask_7_19 = 5'b10000;
localparam output_sel_7_19 = 5'b01000;
localparam input_mask_7_20 = 5'b11000;
localparam output_sel_7_20 = 5'b00100;
localparam input_mask_7_21 = 5'b10100;
localparam output_sel_7_21 = 5'b01000;
localparam input_mask_7_22 = 5'b01000;
localparam output_sel_7_22 = 5'b10000;
localparam input_mask_7_23 = 5'b10000;
localparam output_sel_7_23 = 5'b01000;
localparam input_mask_7_24 = 5'b10000;
localparam output_sel_7_24 = 5'b00000;
localparam input_mask_8_0 = 5'b10000;
localparam output_sel_8_0 = 5'b00000;
localparam input_mask_8_1 = 5'b10000;
localparam output_sel_8_1 = 5'b00000;
localparam input_mask_8_2 = 5'b01000;
localparam output_sel_8_2 = 5'b10000;
localparam input_mask_8_3 = 5'b10000;
localparam output_sel_8_3 = 5'b00000;
localparam input_mask_8_4 = 5'b10000;
localparam output_sel_8_4 = 5'b00001;
localparam input_mask_8_5 = 5'b00110;
localparam output_sel_8_5 = 5'b10000;
localparam input_mask_8_6 = 5'b10000;
localparam output_sel_8_6 = 5'b00100;
localparam input_mask_8_7 = 5'b10000;
localparam output_sel_8_7 = 5'b00100;
localparam input_mask_8_8 = 5'b10000;
localparam output_sel_8_8 = 5'b00001;
localparam input_mask_8_9 = 5'b10010;
localparam output_sel_8_9 = 5'b00100;
localparam input_mask_8_10 = 5'b11000;
localparam output_sel_8_10 = 5'b00100;
localparam input_mask_8_11 = 5'b11000;
localparam output_sel_8_11 = 5'b00100;
localparam input_mask_8_12 = 5'b11000;
localparam output_sel_8_12 = 5'b00100;
localparam input_mask_8_13 = 5'b11000;
localparam output_sel_8_13 = 5'b00100;
localparam input_mask_8_14 = 5'b10000;
localparam output_sel_8_14 = 5'b00100;
localparam input_mask_8_15 = 5'b00100;
localparam output_sel_8_15 = 5'b10000;
localparam input_mask_8_16 = 5'b11000;
localparam output_sel_8_16 = 5'b00100;
localparam input_mask_8_17 = 5'b10100;
localparam output_sel_8_17 = 5'b01000;
localparam input_mask_8_18 = 5'b10000;
localparam output_sel_8_18 = 5'b00100;
localparam input_mask_8_19 = 5'b10000;
localparam output_sel_8_19 = 5'b00100;
localparam input_mask_8_20 = 5'b11000;
localparam output_sel_8_20 = 5'b00100;
localparam input_mask_8_21 = 5'b10100;
localparam output_sel_8_21 = 5'b01000;
localparam input_mask_8_22 = 5'b10000;
localparam output_sel_8_22 = 5'b00100;
localparam input_mask_8_23 = 5'b00100;
localparam output_sel_8_23 = 5'b10000;
localparam input_mask_8_24 = 5'b10000;
localparam output_sel_8_24 = 5'b00000;
localparam input_mask_9_0 = 5'b10000;
localparam output_sel_9_0 = 5'b00000;
localparam input_mask_9_1 = 5'b10000;
localparam output_sel_9_1 = 5'b00000;
localparam input_mask_9_2 = 5'b10000;
localparam output_sel_9_2 = 5'b00000;
localparam input_mask_9_3 = 5'b10000;
localparam output_sel_9_3 = 5'b00000;
localparam input_mask_9_4 = 5'b10000;
localparam output_sel_9_4 = 5'b00001;
localparam input_mask_9_5 = 5'b10010;
localparam output_sel_9_5 = 5'b01000;
localparam input_mask_9_6 = 5'b11000;
localparam output_sel_9_6 = 5'b00001;
localparam input_mask_9_7 = 5'b01010;
localparam output_sel_9_7 = 5'b10000;
localparam input_mask_9_8 = 5'b10000;
localparam output_sel_9_8 = 5'b00001;
localparam input_mask_9_9 = 5'b01010;
localparam output_sel_9_9 = 5'b10000;
localparam input_mask_9_10 = 5'b01000;
localparam output_sel_9_10 = 5'b10000;
localparam input_mask_9_11 = 5'b01000;
localparam output_sel_9_11 = 5'b10000;
localparam input_mask_9_12 = 5'b01000;
localparam output_sel_9_12 = 5'b10000;
localparam input_mask_9_13 = 5'b01000;
localparam output_sel_9_13 = 5'b10000;
localparam input_mask_9_14 = 5'b01000;
localparam output_sel_9_14 = 5'b10000;
localparam input_mask_9_15 = 5'b10000;
localparam output_sel_9_15 = 5'b01000;
localparam input_mask_9_16 = 5'b01000;
localparam output_sel_9_16 = 5'b10000;
localparam input_mask_9_17 = 5'b10000;
localparam output_sel_9_17 = 5'b01000;
localparam input_mask_9_18 = 5'b01000;
localparam output_sel_9_18 = 5'b10000;
localparam input_mask_9_19 = 5'b01000;
localparam output_sel_9_19 = 5'b10000;
localparam input_mask_9_20 = 5'b01000;
localparam output_sel_9_20 = 5'b10000;
localparam input_mask_9_21 = 5'b10000;
localparam output_sel_9_21 = 5'b01000;
localparam input_mask_9_22 = 5'b01000;
localparam output_sel_9_22 = 5'b10000;
localparam input_mask_9_23 = 5'b10000;
localparam output_sel_9_23 = 5'b01000;
localparam input_mask_9_24 = 5'b10000;
localparam output_sel_9_24 = 5'b00000;
`endif
