
`ifndef __NETWORK_CONFIG_SVH_
`define __NETWORK_CONFIG_SVH_
localparam isUBM_list_0_0[`CN] = '{0,0,0,0,0};
localparam isUBM_list_0_1[`CN] = '{0,0,0,0,0};
localparam isUBM_list_0_2[`CN] = '{0,0,0,0,0};
localparam isUBM_list_0_3[`CN] = '{0,0,0,0,0};
localparam isUBM_list_0_4[`CN] = '{0,0,0,0,0};
localparam isUBM_list_0_5[`CN] = '{0,0,0,0,0};
localparam isUBM_list_0_6[`CN] = '{0,0,0,0,0};
localparam isUBM_list_0_7[`CN] = '{0,0,0,0,0};
localparam isUBM_list_1_0[`CN] = '{0,0,0,0,0};
localparam isUBM_list_1_1[`CN] = '{0,0,0,0,0};
localparam isUBM_list_1_2[`CN] = '{0,0,0,0,0};
localparam isUBM_list_1_3[`CN] = '{0,0,0,0,0};
localparam isUBM_list_1_4[`CN] = '{0,0,0,0,0};
localparam isUBM_list_1_5[`CN] = '{0,0,0,0,0};
localparam isUBM_list_1_6[`CN] = '{0,0,0,0,0};
localparam isUBM_list_1_7[`CN] = '{0,0,0,0,0};
localparam isUBM_list_2_0[`CN] = '{0,0,0,0,0};
localparam isUBM_list_2_1[`CN] = '{0,0,0,0,0};
localparam isUBM_list_2_2[`CN] = '{0,0,0,0,0};
localparam isUBM_list_2_3[`CN] = '{0,0,0,0,0};
localparam isUBM_list_2_4[`CN] = '{0,0,0,0,0};
localparam isUBM_list_2_5[`CN] = '{0,0,0,0,0};
localparam isUBM_list_2_6[`CN] = '{0,0,0,0,0};
localparam isUBM_list_2_7[`CN] = '{0,0,0,0,0};
localparam isUBM_list_3_0[`CN] = '{0,0,0,0,0};
localparam isUBM_list_3_1[`CN] = '{0,1,0,0,0};
localparam isUBM_list_3_2[`CN] = '{0,0,0,0,0};
localparam isUBM_list_3_3[`CN] = '{0,0,0,0,0};
localparam isUBM_list_3_4[`CN] = '{1,0,0,0,0};
localparam isUBM_list_3_5[`CN] = '{0,0,0,0,0};
localparam isUBM_list_3_6[`CN] = '{0,0,0,0,0};
localparam isUBM_list_3_7[`CN] = '{0,0,0,0,0};
localparam isUBM_list_4_0[`CN] = '{0,0,0,0,0};
localparam isUBM_list_4_1[`CN] = '{0,0,0,0,0};
localparam isUBM_list_4_2[`CN] = '{0,0,0,0,0};
localparam isUBM_list_4_3[`CN] = '{0,0,0,0,0};
localparam isUBM_list_4_4[`CN] = '{0,0,0,0,0};
localparam isUBM_list_4_5[`CN] = '{0,0,0,0,0};
localparam isUBM_list_4_6[`CN] = '{0,0,0,0,0};
localparam isUBM_list_4_7[`CN] = '{0,0,0,0,0};
localparam isUBM_list_5_0[`CN] = '{0,0,0,0,0};
localparam isUBM_list_5_1[`CN] = '{0,0,0,0,0};
localparam isUBM_list_5_2[`CN] = '{0,0,0,0,0};
localparam isUBM_list_5_3[`CN] = '{0,0,0,0,0};
localparam isUBM_list_5_4[`CN] = '{0,0,0,0,0};
localparam isUBM_list_5_5[`CN] = '{0,0,0,0,0};
localparam isUBM_list_5_6[`CN] = '{0,0,0,0,0};
localparam isUBM_list_5_7[`CN] = '{0,0,0,0,0};
localparam isUBM_list_6_0[`CN] = '{0,0,0,0,0};
localparam isUBM_list_6_1[`CN] = '{0,0,0,0,0};
localparam isUBM_list_6_2[`CN] = '{0,0,0,0,0};
localparam isUBM_list_6_3[`CN] = '{0,0,0,0,0};
localparam isUBM_list_6_4[`CN] = '{0,0,0,0,0};
localparam isUBM_list_6_5[`CN] = '{0,0,0,0,0};
localparam isUBM_list_6_6[`CN] = '{0,0,0,0,0};
localparam isUBM_list_6_7[`CN] = '{0,0,0,0,0};
localparam isFC_list_0_0[`CN] = '{0,0,0,0,0};
localparam isFC_list_0_1[`CN] = '{0,0,0,0,0};
localparam isFC_list_0_2[`CN] = '{0,0,0,0,0};
localparam isFC_list_0_3[`CN] = '{0,0,0,0,0};
localparam isFC_list_0_4[`CN] = '{1,0,0,0,0};
localparam isFC_list_0_5[`CN] = '{0,0,0,0,0};
localparam isFC_list_0_6[`CN] = '{1,0,0,0,0};
localparam isFC_list_0_7[`CN] = '{0,0,0,0,0};
localparam isFC_list_1_0[`CN] = '{0,0,0,0,0};
localparam isFC_list_1_1[`CN] = '{1,0,0,0,0};
localparam isFC_list_1_2[`CN] = '{1,0,0,0,0};
localparam isFC_list_1_3[`CN] = '{0,0,0,0,0};
localparam isFC_list_1_4[`CN] = '{0,0,0,0,0};
localparam isFC_list_1_5[`CN] = '{0,0,0,0,0};
localparam isFC_list_1_6[`CN] = '{0,0,0,0,0};
localparam isFC_list_1_7[`CN] = '{0,0,0,0,0};
localparam isFC_list_2_0[`CN] = '{0,0,0,0,0};
localparam isFC_list_2_1[`CN] = '{0,0,0,0,0};
localparam isFC_list_2_2[`CN] = '{0,0,0,0,0};
localparam isFC_list_2_3[`CN] = '{0,0,0,0,0};
localparam isFC_list_2_4[`CN] = '{0,0,0,0,0};
localparam isFC_list_2_5[`CN] = '{0,0,0,0,0};
localparam isFC_list_2_6[`CN] = '{0,0,0,0,0};
localparam isFC_list_2_7[`CN] = '{0,0,0,0,0};
localparam isFC_list_3_0[`CN] = '{0,0,0,0,0};
localparam isFC_list_3_1[`CN] = '{1,0,0,0,0};
localparam isFC_list_3_2[`CN] = '{0,0,0,0,0};
localparam isFC_list_3_3[`CN] = '{1,0,0,0,0};
localparam isFC_list_3_4[`CN] = '{1,0,0,0,0};
localparam isFC_list_3_5[`CN] = '{0,0,0,0,0};
localparam isFC_list_3_6[`CN] = '{0,0,0,0,0};
localparam isFC_list_3_7[`CN] = '{0,0,0,0,0};
localparam isFC_list_4_0[`CN] = '{1,0,0,0,0};
localparam isFC_list_4_1[`CN] = '{0,0,0,0,0};
localparam isFC_list_4_2[`CN] = '{0,0,0,0,0};
localparam isFC_list_4_3[`CN] = '{0,0,0,0,0};
localparam isFC_list_4_4[`CN] = '{0,0,0,0,0};
localparam isFC_list_4_5[`CN] = '{1,0,0,0,0};
localparam isFC_list_4_6[`CN] = '{0,0,0,0,0};
localparam isFC_list_4_7[`CN] = '{0,0,0,0,0};
localparam isFC_list_5_0[`CN] = '{1,0,0,0,0};
localparam isFC_list_5_1[`CN] = '{0,0,0,0,0};
localparam isFC_list_5_2[`CN] = '{0,0,0,0,0};
localparam isFC_list_5_3[`CN] = '{0,0,0,0,0};
localparam isFC_list_5_4[`CN] = '{0,0,0,0,0};
localparam isFC_list_5_5[`CN] = '{1,0,0,0,0};
localparam isFC_list_5_6[`CN] = '{0,0,0,0,0};
localparam isFC_list_5_7[`CN] = '{0,0,0,0,0};
localparam isFC_list_6_0[`CN] = '{0,0,0,0,0};
localparam isFC_list_6_1[`CN] = '{0,0,0,0,0};
localparam isFC_list_6_2[`CN] = '{0,0,0,0,0};
localparam isFC_list_6_3[`CN] = '{0,0,0,0,0};
localparam isFC_list_6_4[`CN] = '{0,0,0,0,0};
localparam isFC_list_6_5[`CN] = '{0,0,0,0,0};
localparam isFC_list_6_6[`CN] = '{0,0,0,0,0};
localparam isFC_list_6_7[`CN] = '{0,0,0,0,0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_0_0[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_0_1[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_0_2[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_0_3[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_0_4[`CN] = '{56'b00000000000000010000010100100000000000000000000000000000,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_0_5[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_0_6[`CN] = '{56'b10100000110000000000000000000000000000000000000000000000,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_0_7[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_1_0[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_1_1[`CN] = '{56'b00000000000000000000000000000000000110010000000010000000,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_1_2[`CN] = '{56'b00000000000000000000000000011100010000000000000000000000,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_1_3[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_1_4[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_1_5[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_1_6[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_1_7[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_2_0[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_2_1[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_2_2[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_2_3[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_2_4[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_2_5[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_2_6[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_2_7[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_3_0[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_3_1[`CN] = '{56'b00000000000000000000000000000000000001101100000000000000,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_3_2[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_3_3[`CN] = '{56'b00000000000000100000001011000000000000000000000000000000,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_3_4[`CN] = '{56'b00000000000101001100000000000000000000000000000000000000,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_3_5[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_3_6[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_3_7[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_4_0[`CN] = '{56'b00000000000000000000000000000000000000000000000001100000,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_4_1[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_4_2[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_4_3[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_4_4[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_4_5[`CN] = '{56'b01010001001000000000000000000000000000000000000000000000,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_4_6[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_4_7[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_5_0[`CN] = '{56'b00000000000000000000000000000000000000000011000000000000,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_5_1[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_5_2[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_5_3[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_5_4[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_5_5[`CN] = '{56'b00000000000010000011100000000000000000000000000000000000,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_5_6[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_5_7[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_6_0[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_6_1[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_6_2[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_6_3[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_6_4[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_6_5[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_6_6[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_6_7[`CN] = '{56'b0,56'b0,56'b0,56'b0,56'b0};
localparam int FCpl_list_0_0[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_0_1[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_0_2[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_0_3[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_0_4[`CN] = '{`PKT_LEN,0,0,0,0};
localparam int FCpl_list_0_5[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_0_6[`CN] = '{`PKT_LEN,0,0,0,0};
localparam int FCpl_list_0_7[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_1_0[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_1_1[`CN] = '{`PKT_LEN,0,0,0,0};
localparam int FCpl_list_1_2[`CN] = '{`PKT_LEN,0,0,0,0};
localparam int FCpl_list_1_3[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_1_4[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_1_5[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_1_6[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_1_7[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_2_0[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_2_1[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_2_2[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_2_3[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_2_4[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_2_5[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_2_6[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_2_7[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_3_0[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_3_1[`CN] = '{`PKT_LEN,0,0,0,0};
localparam int FCpl_list_3_2[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_3_3[`CN] = '{`PKT_LEN,0,0,0,0};
localparam int FCpl_list_3_4[`CN] = '{`PKT_LEN,0,0,0,0};
localparam int FCpl_list_3_5[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_3_6[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_3_7[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_4_0[`CN] = '{`PKT_LEN,0,0,0,0};
localparam int FCpl_list_4_1[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_4_2[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_4_3[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_4_4[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_4_5[`CN] = '{`PKT_LEN,0,0,0,0};
localparam int FCpl_list_4_6[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_4_7[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_5_0[`CN] = '{`PKT_LEN,0,0,0,0};
localparam int FCpl_list_5_1[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_5_2[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_5_3[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_5_4[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_5_5[`CN] = '{`PKT_LEN,0,0,0,0};
localparam int FCpl_list_5_6[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_5_7[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_6_0[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_6_1[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_6_2[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_6_3[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_6_4[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_6_5[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_6_6[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_6_7[`CN] = '{0,0,0,0,0};
localparam string rt_file_list_0_0[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_0_0_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_0_0_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_0_0_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_0_0_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_0_0_4"};
localparam string rt_file_list_0_1[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_0_1_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_0_1_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_0_1_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_0_1_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_0_1_4"};
localparam string rt_file_list_0_2[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_0_2_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_0_2_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_0_2_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_0_2_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_0_2_4"};
localparam string rt_file_list_0_3[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_0_3_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_0_3_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_0_3_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_0_3_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_0_3_4"};
localparam string rt_file_list_0_4[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_0_4_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_0_4_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_0_4_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_0_4_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_0_4_4"};
localparam string rt_file_list_0_5[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_0_5_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_0_5_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_0_5_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_0_5_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_0_5_4"};
localparam string rt_file_list_0_6[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_0_6_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_0_6_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_0_6_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_0_6_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_0_6_4"};
localparam string rt_file_list_0_7[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_0_7_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_0_7_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_0_7_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_0_7_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_0_7_4"};
localparam string rt_file_list_1_0[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_1_0_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_1_0_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_1_0_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_1_0_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_1_0_4"};
localparam string rt_file_list_1_1[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_1_1_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_1_1_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_1_1_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_1_1_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_1_1_4"};
localparam string rt_file_list_1_2[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_1_2_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_1_2_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_1_2_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_1_2_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_1_2_4"};
localparam string rt_file_list_1_3[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_1_3_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_1_3_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_1_3_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_1_3_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_1_3_4"};
localparam string rt_file_list_1_4[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_1_4_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_1_4_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_1_4_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_1_4_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_1_4_4"};
localparam string rt_file_list_1_5[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_1_5_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_1_5_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_1_5_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_1_5_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_1_5_4"};
localparam string rt_file_list_1_6[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_1_6_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_1_6_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_1_6_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_1_6_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_1_6_4"};
localparam string rt_file_list_1_7[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_1_7_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_1_7_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_1_7_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_1_7_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_1_7_4"};
localparam string rt_file_list_2_0[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_2_0_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_2_0_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_2_0_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_2_0_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_2_0_4"};
localparam string rt_file_list_2_1[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_2_1_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_2_1_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_2_1_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_2_1_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_2_1_4"};
localparam string rt_file_list_2_2[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_2_2_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_2_2_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_2_2_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_2_2_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_2_2_4"};
localparam string rt_file_list_2_3[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_2_3_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_2_3_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_2_3_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_2_3_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_2_3_4"};
localparam string rt_file_list_2_4[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_2_4_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_2_4_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_2_4_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_2_4_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_2_4_4"};
localparam string rt_file_list_2_5[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_2_5_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_2_5_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_2_5_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_2_5_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_2_5_4"};
localparam string rt_file_list_2_6[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_2_6_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_2_6_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_2_6_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_2_6_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_2_6_4"};
localparam string rt_file_list_2_7[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_2_7_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_2_7_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_2_7_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_2_7_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_2_7_4"};
localparam string rt_file_list_3_0[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_3_0_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_3_0_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_3_0_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_3_0_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_3_0_4"};
localparam string rt_file_list_3_1[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_3_1_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_3_1_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_3_1_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_3_1_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_3_1_4"};
localparam string rt_file_list_3_2[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_3_2_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_3_2_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_3_2_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_3_2_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_3_2_4"};
localparam string rt_file_list_3_3[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_3_3_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_3_3_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_3_3_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_3_3_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_3_3_4"};
localparam string rt_file_list_3_4[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_3_4_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_3_4_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_3_4_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_3_4_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_3_4_4"};
localparam string rt_file_list_3_5[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_3_5_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_3_5_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_3_5_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_3_5_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_3_5_4"};
localparam string rt_file_list_3_6[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_3_6_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_3_6_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_3_6_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_3_6_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_3_6_4"};
localparam string rt_file_list_3_7[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_3_7_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_3_7_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_3_7_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_3_7_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_3_7_4"};
localparam string rt_file_list_4_0[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_4_0_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_4_0_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_4_0_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_4_0_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_4_0_4"};
localparam string rt_file_list_4_1[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_4_1_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_4_1_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_4_1_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_4_1_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_4_1_4"};
localparam string rt_file_list_4_2[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_4_2_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_4_2_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_4_2_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_4_2_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_4_2_4"};
localparam string rt_file_list_4_3[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_4_3_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_4_3_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_4_3_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_4_3_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_4_3_4"};
localparam string rt_file_list_4_4[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_4_4_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_4_4_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_4_4_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_4_4_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_4_4_4"};
localparam string rt_file_list_4_5[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_4_5_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_4_5_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_4_5_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_4_5_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_4_5_4"};
localparam string rt_file_list_4_6[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_4_6_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_4_6_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_4_6_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_4_6_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_4_6_4"};
localparam string rt_file_list_4_7[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_4_7_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_4_7_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_4_7_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_4_7_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_4_7_4"};
localparam string rt_file_list_5_0[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_5_0_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_5_0_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_5_0_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_5_0_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_5_0_4"};
localparam string rt_file_list_5_1[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_5_1_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_5_1_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_5_1_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_5_1_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_5_1_4"};
localparam string rt_file_list_5_2[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_5_2_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_5_2_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_5_2_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_5_2_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_5_2_4"};
localparam string rt_file_list_5_3[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_5_3_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_5_3_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_5_3_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_5_3_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_5_3_4"};
localparam string rt_file_list_5_4[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_5_4_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_5_4_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_5_4_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_5_4_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_5_4_4"};
localparam string rt_file_list_5_5[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_5_5_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_5_5_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_5_5_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_5_5_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_5_5_4"};
localparam string rt_file_list_5_6[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_5_6_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_5_6_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_5_6_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_5_6_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_5_6_4"};
localparam string rt_file_list_5_7[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_5_7_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_5_7_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_5_7_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_5_7_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_5_7_4"};
localparam string rt_file_list_6_0[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_6_0_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_6_0_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_6_0_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_6_0_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_6_0_4"};
localparam string rt_file_list_6_1[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_6_1_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_6_1_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_6_1_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_6_1_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_6_1_4"};
localparam string rt_file_list_6_2[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_6_2_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_6_2_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_6_2_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_6_2_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_6_2_4"};
localparam string rt_file_list_6_3[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_6_3_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_6_3_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_6_3_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_6_3_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_6_3_4"};
localparam string rt_file_list_6_4[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_6_4_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_6_4_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_6_4_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_6_4_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_6_4_4"};
localparam string rt_file_list_6_5[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_6_5_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_6_5_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_6_5_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_6_5_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_6_5_4"};
localparam string rt_file_list_6_6[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_6_6_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_6_6_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_6_6_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_6_6_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_6_6_4"};
localparam string rt_file_list_6_7[`CN] = '{"/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_6_7_0","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_6_7_1","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_6_7_2","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_6_7_3","/mnt/c/git/nvcim-comm/network/srcs/config/cast_rt_6_7_4"};


localparam input_mask_0_0 = 5'b00000;
localparam output_sel_0_0 = 5'b00001;
localparam input_mask_0_1 = 5'b00001;
localparam output_sel_0_1 = 5'b10000;
localparam input_mask_0_2 = 5'b01001;
localparam output_sel_0_2 = 5'b00100;
localparam input_mask_0_3 = 5'b00101;
localparam output_sel_0_3 = 5'b10000;
localparam input_mask_0_4 = 5'b01000;
localparam output_sel_0_4 = 5'b00001;
localparam input_mask_0_5 = 5'b00001;
localparam output_sel_0_5 = 5'b10000;
localparam input_mask_0_6 = 5'b01100;
localparam output_sel_0_6 = 5'b00001;
localparam input_mask_0_7 = 5'b00000;
localparam output_sel_0_7 = 5'b00001;
localparam input_mask_1_0 = 5'b00000;
localparam output_sel_1_0 = 5'b00001;
localparam input_mask_1_1 = 5'b00100;
localparam output_sel_1_1 = 5'b00001;
localparam input_mask_1_2 = 5'b00110;
localparam output_sel_1_2 = 5'b00001;
localparam input_mask_1_3 = 5'b00101;
localparam output_sel_1_3 = 5'b00010;
localparam input_mask_1_4 = 5'b00001;
localparam output_sel_1_4 = 5'b00100;
localparam input_mask_1_5 = 5'b00001;
localparam output_sel_1_5 = 5'b00100;
localparam input_mask_1_6 = 5'b00101;
localparam output_sel_1_6 = 5'b00010;
localparam input_mask_1_7 = 5'b00000;
localparam output_sel_1_7 = 5'b00001;
localparam input_mask_2_0 = 5'b00000;
localparam output_sel_2_0 = 5'b00001;
localparam input_mask_2_1 = 5'b00001;
localparam output_sel_2_1 = 5'b00010;
localparam input_mask_2_2 = 5'b00001;
localparam output_sel_2_2 = 5'b00010;
localparam input_mask_2_3 = 5'b00001;
localparam output_sel_2_3 = 5'b00010;
localparam input_mask_2_4 = 5'b00011;
localparam output_sel_2_4 = 5'b00100;
localparam input_mask_2_5 = 5'b00011;
localparam output_sel_2_5 = 5'b00100;
localparam input_mask_2_6 = 5'b00001;
localparam output_sel_2_6 = 5'b00010;
localparam input_mask_2_7 = 5'b00000;
localparam output_sel_2_7 = 5'b00001;
localparam input_mask_3_0 = 5'b00000;
localparam output_sel_3_0 = 5'b00001;
localparam input_mask_3_1 = 5'b00100;
localparam output_sel_3_1 = 5'b00001;
localparam input_mask_3_2 = 5'b00001;
localparam output_sel_3_2 = 5'b00100;
localparam input_mask_3_3 = 5'b00100;
localparam output_sel_3_3 = 5'b00001;
localparam input_mask_3_4 = 5'b00110;
localparam output_sel_3_4 = 5'b00001;
localparam input_mask_3_5 = 5'b00011;
localparam output_sel_3_5 = 5'b00100;
localparam input_mask_3_6 = 5'b00001;
localparam output_sel_3_6 = 5'b00100;
localparam input_mask_3_7 = 5'b00001;
localparam output_sel_3_7 = 5'b00100;
localparam input_mask_4_0 = 5'b00000;
localparam output_sel_4_0 = 5'b00001;
localparam input_mask_4_1 = 5'b00001;
localparam output_sel_4_1 = 5'b00010;
localparam input_mask_4_2 = 5'b00011;
localparam output_sel_4_2 = 5'b00100;
localparam input_mask_4_3 = 5'b00101;
localparam output_sel_4_3 = 5'b00010;
localparam input_mask_4_4 = 5'b00001;
localparam output_sel_4_4 = 5'b00010;
localparam input_mask_4_5 = 5'b00010;
localparam output_sel_4_5 = 5'b00001;
localparam input_mask_4_6 = 5'b00011;
localparam output_sel_4_6 = 5'b00100;
localparam input_mask_4_7 = 5'b00110;
localparam output_sel_4_7 = 5'b00001;
localparam input_mask_5_0 = 5'b00100;
localparam output_sel_5_0 = 5'b00001;
localparam input_mask_5_1 = 5'b00100;
localparam output_sel_5_1 = 5'b00001;
localparam input_mask_5_2 = 5'b00011;
localparam output_sel_5_2 = 5'b00100;
localparam input_mask_5_3 = 5'b00101;
localparam output_sel_5_3 = 5'b00010;
localparam input_mask_5_4 = 5'b00001;
localparam output_sel_5_4 = 5'b10000;
localparam input_mask_5_5 = 5'b01100;
localparam output_sel_5_5 = 5'b00001;
localparam input_mask_5_6 = 5'b00011;
localparam output_sel_5_6 = 5'b00100;
localparam input_mask_5_7 = 5'b00101;
localparam output_sel_5_7 = 5'b00010;
localparam input_mask_6_0 = 5'b00001;
localparam output_sel_6_0 = 5'b00010;
localparam input_mask_6_1 = 5'b00001;
localparam output_sel_6_1 = 5'b00010;
localparam input_mask_6_2 = 5'b00010;
localparam output_sel_6_2 = 5'b00001;
localparam input_mask_6_3 = 5'b00001;
localparam output_sel_6_3 = 5'b00010;
localparam input_mask_6_4 = 5'b00001;
localparam output_sel_6_4 = 5'b10000;
localparam input_mask_6_5 = 5'b01001;
localparam output_sel_6_5 = 5'b00010;
localparam input_mask_6_6 = 5'b00010;
localparam output_sel_6_6 = 5'b00001;
localparam input_mask_6_7 = 5'b00001;
localparam output_sel_6_7 = 5'b00010;


localparam isCaster_0_0 = 1;
localparam stream_id_0_0 = 1;
localparam isCaster_0_1 = 0;
localparam stream_id_0_1 = 0;
localparam isCaster_0_2 = 0;
localparam stream_id_0_2 = 0;
localparam isCaster_0_3 = 0;
localparam stream_id_0_3 = 0;
localparam isCaster_0_4 = 1;
localparam stream_id_0_4 = 13;
localparam isCaster_0_5 = 0;
localparam stream_id_0_5 = 0;
localparam isCaster_0_6 = 1;
localparam stream_id_0_6 = 17;
localparam isCaster_0_7 = 0;
localparam stream_id_0_7 = 0;
localparam isCaster_1_0 = 1;
localparam stream_id_1_0 = 2;
localparam isCaster_1_1 = 1;
localparam stream_id_1_1 = 9;
localparam isCaster_1_2 = 1;
localparam stream_id_1_2 = 10;
localparam isCaster_1_3 = 0;
localparam stream_id_1_3 = 0;
localparam isCaster_1_4 = 0;
localparam stream_id_1_4 = 0;
localparam isCaster_1_5 = 0;
localparam stream_id_1_5 = 0;
localparam isCaster_1_6 = 0;
localparam stream_id_1_6 = 0;
localparam isCaster_1_7 = 0;
localparam stream_id_1_7 = 0;
localparam isCaster_2_0 = 1;
localparam stream_id_2_0 = 3;
localparam isCaster_2_1 = 0;
localparam stream_id_2_1 = 0;
localparam isCaster_2_2 = 0;
localparam stream_id_2_2 = 0;
localparam isCaster_2_3 = 0;
localparam stream_id_2_3 = 0;
localparam isCaster_2_4 = 0;
localparam stream_id_2_4 = 0;
localparam isCaster_2_5 = 0;
localparam stream_id_2_5 = 0;
localparam isCaster_2_6 = 0;
localparam stream_id_2_6 = 0;
localparam isCaster_2_7 = 0;
localparam stream_id_2_7 = 0;
localparam isCaster_3_0 = 1;
localparam stream_id_3_0 = 4;
localparam isCaster_3_1 = 1;
localparam stream_id_3_1 = 8;
localparam isCaster_3_2 = 0;
localparam stream_id_3_2 = 0;
localparam isCaster_3_3 = 1;
localparam stream_id_3_3 = 12;
localparam isCaster_3_4 = 1;
localparam stream_id_3_4 = 14;
localparam isCaster_3_5 = 0;
localparam stream_id_3_5 = 0;
localparam isCaster_3_6 = 0;
localparam stream_id_3_6 = 0;
localparam isCaster_3_7 = 0;
localparam stream_id_3_7 = 0;
localparam isCaster_4_0 = 1;
localparam stream_id_4_0 = 5;
localparam isCaster_4_1 = 0;
localparam stream_id_4_1 = 0;
localparam isCaster_4_2 = 0;
localparam stream_id_4_2 = 0;
localparam isCaster_4_3 = 0;
localparam stream_id_4_3 = 0;
localparam isCaster_4_4 = 0;
localparam stream_id_4_4 = 0;
localparam isCaster_4_5 = 1;
localparam stream_id_4_5 = 16;
localparam isCaster_4_6 = 0;
localparam stream_id_4_6 = 0;
localparam isCaster_4_7 = 1;
localparam stream_id_4_7 = 1022;
localparam isCaster_5_0 = 1;
localparam stream_id_5_0 = 6;
localparam isCaster_5_1 = 1;
localparam stream_id_5_1 = 7;
localparam isCaster_5_2 = 0;
localparam stream_id_5_2 = 0;
localparam isCaster_5_3 = 0;
localparam stream_id_5_3 = 0;
localparam isCaster_5_4 = 0;
localparam stream_id_5_4 = 0;
localparam isCaster_5_5 = 1;
localparam stream_id_5_5 = 15;
localparam isCaster_5_6 = 0;
localparam stream_id_5_6 = 0;
localparam isCaster_5_7 = 0;
localparam stream_id_5_7 = 0;
localparam isCaster_6_0 = 0;
localparam stream_id_6_0 = 0;
localparam isCaster_6_1 = 0;
localparam stream_id_6_1 = 0;
localparam isCaster_6_2 = 1;
localparam stream_id_6_2 = 11;
localparam isCaster_6_3 = 0;
localparam stream_id_6_3 = 0;
localparam isCaster_6_4 = 0;
localparam stream_id_6_4 = 0;
localparam isCaster_6_5 = 0;
localparam stream_id_6_5 = 0;
localparam isCaster_6_6 = 1;
localparam stream_id_6_6 = 1022;
localparam isCaster_6_7 = 0;
localparam stream_id_6_7 = 0;

`endif
        
