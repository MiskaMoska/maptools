
//Cast Network
//Width: 5
//Height:10
`include "params.svh"
`include "cast_network_config.svh"

module cast_network(
    input       wire                            clk,
    input       wire                            rstn,

    //router local ports
    input       wire        [`DW-1:0]           data_i[`NOC_WIDTH][`NOC_HEIGHT],
    input       wire                            valid_i[`NOC_WIDTH][`NOC_HEIGHT],
    output      wire                            ready_o[`NOC_WIDTH][`NOC_HEIGHT],

    output      wire        [`DW-1:0]           data_o[`NOC_WIDTH][`NOC_HEIGHT],
    output      wire                            valid_o[`NOC_WIDTH][`NOC_HEIGHT],
    input       wire                            ready_i[`NOC_WIDTH][`NOC_HEIGHT],

    input       wire        [`DW-1:0]           data_i_stab,
    input       wire                            valid_i_stab,
    output      wire                            ready_o_stab,

    output      wire        [`DW-1:0]           data_o_flee0,
    output      wire                            valid_o_flee0,
    input       wire                            ready_i_flee0,

    output      wire        [`DW-1:0]           data_o_flee1,
    output      wire                            valid_o_flee1,
    input       wire                            ready_i_flee1,

    //credit update signal input
    input       wire                            credit_upd[`NOC_WIDTH][`NOC_HEIGHT]

);

//horizontal signals
wire    [`DW-1:0]   data_0_to_1,	data_1_to_0;
wire                valid_0_to_1,	valid_1_to_0;
wire                ready_0_to_1,	ready_1_to_0;
wire    [`DW-1:0]   data_1_to_2,	data_2_to_1;
wire                valid_1_to_2,	valid_2_to_1;
wire                ready_1_to_2,	ready_2_to_1;
wire    [`DW-1:0]   data_2_to_3,	data_3_to_2;
wire                valid_2_to_3,	valid_3_to_2;
wire                ready_2_to_3,	ready_3_to_2;
wire    [`DW-1:0]   data_3_to_4,	data_4_to_3;
wire                valid_3_to_4,	valid_4_to_3;
wire                ready_3_to_4,	ready_4_to_3;
wire    [`DW-1:0]   data_5_to_6,	data_6_to_5;
wire                valid_5_to_6,	valid_6_to_5;
wire                ready_5_to_6,	ready_6_to_5;
wire    [`DW-1:0]   data_6_to_7,	data_7_to_6;
wire                valid_6_to_7,	valid_7_to_6;
wire                ready_6_to_7,	ready_7_to_6;
wire    [`DW-1:0]   data_7_to_8,	data_8_to_7;
wire                valid_7_to_8,	valid_8_to_7;
wire                ready_7_to_8,	ready_8_to_7;
wire    [`DW-1:0]   data_8_to_9,	data_9_to_8;
wire                valid_8_to_9,	valid_9_to_8;
wire                ready_8_to_9,	ready_9_to_8;
wire    [`DW-1:0]   data_10_to_11,	data_11_to_10;
wire                valid_10_to_11,	valid_11_to_10;
wire                ready_10_to_11,	ready_11_to_10;
wire    [`DW-1:0]   data_11_to_12,	data_12_to_11;
wire                valid_11_to_12,	valid_12_to_11;
wire                ready_11_to_12,	ready_12_to_11;
wire    [`DW-1:0]   data_12_to_13,	data_13_to_12;
wire                valid_12_to_13,	valid_13_to_12;
wire                ready_12_to_13,	ready_13_to_12;
wire    [`DW-1:0]   data_13_to_14,	data_14_to_13;
wire                valid_13_to_14,	valid_14_to_13;
wire                ready_13_to_14,	ready_14_to_13;
wire    [`DW-1:0]   data_15_to_16,	data_16_to_15;
wire                valid_15_to_16,	valid_16_to_15;
wire                ready_15_to_16,	ready_16_to_15;
wire    [`DW-1:0]   data_16_to_17,	data_17_to_16;
wire                valid_16_to_17,	valid_17_to_16;
wire                ready_16_to_17,	ready_17_to_16;
wire    [`DW-1:0]   data_17_to_18,	data_18_to_17;
wire                valid_17_to_18,	valid_18_to_17;
wire                ready_17_to_18,	ready_18_to_17;
wire    [`DW-1:0]   data_18_to_19,	data_19_to_18;
wire                valid_18_to_19,	valid_19_to_18;
wire                ready_18_to_19,	ready_19_to_18;
wire    [`DW-1:0]   data_20_to_21,	data_21_to_20;
wire                valid_20_to_21,	valid_21_to_20;
wire                ready_20_to_21,	ready_21_to_20;
wire    [`DW-1:0]   data_21_to_22,	data_22_to_21;
wire                valid_21_to_22,	valid_22_to_21;
wire                ready_21_to_22,	ready_22_to_21;
wire    [`DW-1:0]   data_22_to_23,	data_23_to_22;
wire                valid_22_to_23,	valid_23_to_22;
wire                ready_22_to_23,	ready_23_to_22;
wire    [`DW-1:0]   data_23_to_24,	data_24_to_23;
wire                valid_23_to_24,	valid_24_to_23;
wire                ready_23_to_24,	ready_24_to_23;
wire    [`DW-1:0]   data_25_to_26,	data_26_to_25;
wire                valid_25_to_26,	valid_26_to_25;
wire                ready_25_to_26,	ready_26_to_25;
wire    [`DW-1:0]   data_26_to_27,	data_27_to_26;
wire                valid_26_to_27,	valid_27_to_26;
wire                ready_26_to_27,	ready_27_to_26;
wire    [`DW-1:0]   data_27_to_28,	data_28_to_27;
wire                valid_27_to_28,	valid_28_to_27;
wire                ready_27_to_28,	ready_28_to_27;
wire    [`DW-1:0]   data_28_to_29,	data_29_to_28;
wire                valid_28_to_29,	valid_29_to_28;
wire                ready_28_to_29,	ready_29_to_28;
wire    [`DW-1:0]   data_30_to_31,	data_31_to_30;
wire                valid_30_to_31,	valid_31_to_30;
wire                ready_30_to_31,	ready_31_to_30;
wire    [`DW-1:0]   data_31_to_32,	data_32_to_31;
wire                valid_31_to_32,	valid_32_to_31;
wire                ready_31_to_32,	ready_32_to_31;
wire    [`DW-1:0]   data_32_to_33,	data_33_to_32;
wire                valid_32_to_33,	valid_33_to_32;
wire                ready_32_to_33,	ready_33_to_32;
wire    [`DW-1:0]   data_33_to_34,	data_34_to_33;
wire                valid_33_to_34,	valid_34_to_33;
wire                ready_33_to_34,	ready_34_to_33;
wire    [`DW-1:0]   data_35_to_36,	data_36_to_35;
wire                valid_35_to_36,	valid_36_to_35;
wire                ready_35_to_36,	ready_36_to_35;
wire    [`DW-1:0]   data_36_to_37,	data_37_to_36;
wire                valid_36_to_37,	valid_37_to_36;
wire                ready_36_to_37,	ready_37_to_36;
wire    [`DW-1:0]   data_37_to_38,	data_38_to_37;
wire                valid_37_to_38,	valid_38_to_37;
wire                ready_37_to_38,	ready_38_to_37;
wire    [`DW-1:0]   data_38_to_39,	data_39_to_38;
wire                valid_38_to_39,	valid_39_to_38;
wire                ready_38_to_39,	ready_39_to_38;
wire    [`DW-1:0]   data_40_to_41,	data_41_to_40;
wire                valid_40_to_41,	valid_41_to_40;
wire                ready_40_to_41,	ready_41_to_40;
wire    [`DW-1:0]   data_41_to_42,	data_42_to_41;
wire                valid_41_to_42,	valid_42_to_41;
wire                ready_41_to_42,	ready_42_to_41;
wire    [`DW-1:0]   data_42_to_43,	data_43_to_42;
wire                valid_42_to_43,	valid_43_to_42;
wire                ready_42_to_43,	ready_43_to_42;
wire    [`DW-1:0]   data_43_to_44,	data_44_to_43;
wire                valid_43_to_44,	valid_44_to_43;
wire                ready_43_to_44,	ready_44_to_43;
wire    [`DW-1:0]   data_45_to_46,	data_46_to_45;
wire                valid_45_to_46,	valid_46_to_45;
wire                ready_45_to_46,	ready_46_to_45;
wire    [`DW-1:0]   data_46_to_47,	data_47_to_46;
wire                valid_46_to_47,	valid_47_to_46;
wire                ready_46_to_47,	ready_47_to_46;
wire    [`DW-1:0]   data_47_to_48,	data_48_to_47;
wire                valid_47_to_48,	valid_48_to_47;
wire                ready_47_to_48,	ready_48_to_47;
wire    [`DW-1:0]   data_48_to_49,	data_49_to_48;
wire                valid_48_to_49,	valid_49_to_48;
wire                ready_48_to_49,	ready_49_to_48;

//vertical signals
wire    [`DW-1:0]   data_0_to_5_v0,	data_0_to_5_v1;
wire                valid_0_to_5_v0,	valid_0_to_5_v1;
wire                ready_5_to_0_v0,	ready_5_to_0_v1;
wire    [`DW-1:0]   data_5_to_10_v0,	data_5_to_10_v1;
wire                valid_5_to_10_v0,	valid_5_to_10_v1;
wire                ready_10_to_5_v0,	ready_10_to_5_v1;
wire    [`DW-1:0]   data_10_to_15_v0,	data_10_to_15_v1;
wire                valid_10_to_15_v0,	valid_10_to_15_v1;
wire                ready_15_to_10_v0,	ready_15_to_10_v1;
wire    [`DW-1:0]   data_15_to_20_v0,	data_15_to_20_v1;
wire                valid_15_to_20_v0,	valid_15_to_20_v1;
wire                ready_20_to_15_v0,	ready_20_to_15_v1;
wire    [`DW-1:0]   data_20_to_25_v0,	data_20_to_25_v1;
wire                valid_20_to_25_v0,	valid_20_to_25_v1;
wire                ready_25_to_20_v0,	ready_25_to_20_v1;
wire    [`DW-1:0]   data_25_to_30_v0,	data_25_to_30_v1;
wire                valid_25_to_30_v0,	valid_25_to_30_v1;
wire                ready_30_to_25_v0,	ready_30_to_25_v1;
wire    [`DW-1:0]   data_30_to_35_v0,	data_30_to_35_v1;
wire                valid_30_to_35_v0,	valid_30_to_35_v1;
wire                ready_35_to_30_v0,	ready_35_to_30_v1;
wire    [`DW-1:0]   data_35_to_40_v0,	data_35_to_40_v1;
wire                valid_35_to_40_v0,	valid_35_to_40_v1;
wire                ready_40_to_35_v0,	ready_40_to_35_v1;
wire    [`DW-1:0]   data_40_to_45_v0,	data_40_to_45_v1;
wire                valid_40_to_45_v0,	valid_40_to_45_v1;
wire                ready_45_to_40_v0,	ready_45_to_40_v1;
wire    [`DW-1:0]   data_1_to_6_v0,	data_1_to_6_v1;
wire                valid_1_to_6_v0,	valid_1_to_6_v1;
wire                ready_6_to_1_v0,	ready_6_to_1_v1;
wire    [`DW-1:0]   data_6_to_11_v0,	data_6_to_11_v1;
wire                valid_6_to_11_v0,	valid_6_to_11_v1;
wire                ready_11_to_6_v0,	ready_11_to_6_v1;
wire    [`DW-1:0]   data_11_to_16_v0,	data_11_to_16_v1;
wire                valid_11_to_16_v0,	valid_11_to_16_v1;
wire                ready_16_to_11_v0,	ready_16_to_11_v1;
wire    [`DW-1:0]   data_16_to_21_v0,	data_16_to_21_v1;
wire                valid_16_to_21_v0,	valid_16_to_21_v1;
wire                ready_21_to_16_v0,	ready_21_to_16_v1;
wire    [`DW-1:0]   data_21_to_26_v0,	data_21_to_26_v1;
wire                valid_21_to_26_v0,	valid_21_to_26_v1;
wire                ready_26_to_21_v0,	ready_26_to_21_v1;
wire    [`DW-1:0]   data_26_to_31_v0,	data_26_to_31_v1;
wire                valid_26_to_31_v0,	valid_26_to_31_v1;
wire                ready_31_to_26_v0,	ready_31_to_26_v1;
wire    [`DW-1:0]   data_31_to_36_v0,	data_31_to_36_v1;
wire                valid_31_to_36_v0,	valid_31_to_36_v1;
wire                ready_36_to_31_v0,	ready_36_to_31_v1;
wire    [`DW-1:0]   data_36_to_41_v0,	data_36_to_41_v1;
wire                valid_36_to_41_v0,	valid_36_to_41_v1;
wire                ready_41_to_36_v0,	ready_41_to_36_v1;
wire    [`DW-1:0]   data_41_to_46_v0,	data_41_to_46_v1;
wire                valid_41_to_46_v0,	valid_41_to_46_v1;
wire                ready_46_to_41_v0,	ready_46_to_41_v1;
wire    [`DW-1:0]   data_2_to_7_v0,	data_2_to_7_v1;
wire                valid_2_to_7_v0,	valid_2_to_7_v1;
wire                ready_7_to_2_v0,	ready_7_to_2_v1;
wire    [`DW-1:0]   data_7_to_12_v0,	data_7_to_12_v1;
wire                valid_7_to_12_v0,	valid_7_to_12_v1;
wire                ready_12_to_7_v0,	ready_12_to_7_v1;
wire    [`DW-1:0]   data_12_to_17_v0,	data_12_to_17_v1;
wire                valid_12_to_17_v0,	valid_12_to_17_v1;
wire                ready_17_to_12_v0,	ready_17_to_12_v1;
wire    [`DW-1:0]   data_17_to_22_v0,	data_17_to_22_v1;
wire                valid_17_to_22_v0,	valid_17_to_22_v1;
wire                ready_22_to_17_v0,	ready_22_to_17_v1;
wire    [`DW-1:0]   data_22_to_27_v0,	data_22_to_27_v1;
wire                valid_22_to_27_v0,	valid_22_to_27_v1;
wire                ready_27_to_22_v0,	ready_27_to_22_v1;
wire    [`DW-1:0]   data_27_to_32_v0,	data_27_to_32_v1;
wire                valid_27_to_32_v0,	valid_27_to_32_v1;
wire                ready_32_to_27_v0,	ready_32_to_27_v1;
wire    [`DW-1:0]   data_32_to_37_v0,	data_32_to_37_v1;
wire                valid_32_to_37_v0,	valid_32_to_37_v1;
wire                ready_37_to_32_v0,	ready_37_to_32_v1;
wire    [`DW-1:0]   data_37_to_42_v0,	data_37_to_42_v1;
wire                valid_37_to_42_v0,	valid_37_to_42_v1;
wire                ready_42_to_37_v0,	ready_42_to_37_v1;
wire    [`DW-1:0]   data_42_to_47_v0,	data_42_to_47_v1;
wire                valid_42_to_47_v0,	valid_42_to_47_v1;
wire                ready_47_to_42_v0,	ready_47_to_42_v1;
wire    [`DW-1:0]   data_3_to_8_v0,	data_3_to_8_v1;
wire                valid_3_to_8_v0,	valid_3_to_8_v1;
wire                ready_8_to_3_v0,	ready_8_to_3_v1;
wire    [`DW-1:0]   data_8_to_13_v0,	data_8_to_13_v1;
wire                valid_8_to_13_v0,	valid_8_to_13_v1;
wire                ready_13_to_8_v0,	ready_13_to_8_v1;
wire    [`DW-1:0]   data_13_to_18_v0,	data_13_to_18_v1;
wire                valid_13_to_18_v0,	valid_13_to_18_v1;
wire                ready_18_to_13_v0,	ready_18_to_13_v1;
wire    [`DW-1:0]   data_18_to_23_v0,	data_18_to_23_v1;
wire                valid_18_to_23_v0,	valid_18_to_23_v1;
wire                ready_23_to_18_v0,	ready_23_to_18_v1;
wire    [`DW-1:0]   data_23_to_28_v0,	data_23_to_28_v1;
wire                valid_23_to_28_v0,	valid_23_to_28_v1;
wire                ready_28_to_23_v0,	ready_28_to_23_v1;
wire    [`DW-1:0]   data_28_to_33_v0,	data_28_to_33_v1;
wire                valid_28_to_33_v0,	valid_28_to_33_v1;
wire                ready_33_to_28_v0,	ready_33_to_28_v1;
wire    [`DW-1:0]   data_33_to_38_v0,	data_33_to_38_v1;
wire                valid_33_to_38_v0,	valid_33_to_38_v1;
wire                ready_38_to_33_v0,	ready_38_to_33_v1;
wire    [`DW-1:0]   data_38_to_43_v0,	data_38_to_43_v1;
wire                valid_38_to_43_v0,	valid_38_to_43_v1;
wire                ready_43_to_38_v0,	ready_43_to_38_v1;
wire    [`DW-1:0]   data_43_to_48_v0,	data_43_to_48_v1;
wire                valid_43_to_48_v0,	valid_43_to_48_v1;
wire                ready_48_to_43_v0,	ready_48_to_43_v1;
wire    [`DW-1:0]   data_4_to_9_v0,	data_4_to_9_v1;
wire                valid_4_to_9_v0,	valid_4_to_9_v1;
wire                ready_9_to_4_v0,	ready_9_to_4_v1;
wire    [`DW-1:0]   data_9_to_14_v0,	data_9_to_14_v1;
wire                valid_9_to_14_v0,	valid_9_to_14_v1;
wire                ready_14_to_9_v0,	ready_14_to_9_v1;
wire    [`DW-1:0]   data_14_to_19_v0,	data_14_to_19_v1;
wire                valid_14_to_19_v0,	valid_14_to_19_v1;
wire                ready_19_to_14_v0,	ready_19_to_14_v1;
wire    [`DW-1:0]   data_19_to_24_v0,	data_19_to_24_v1;
wire                valid_19_to_24_v0,	valid_19_to_24_v1;
wire                ready_24_to_19_v0,	ready_24_to_19_v1;
wire    [`DW-1:0]   data_24_to_29_v0,	data_24_to_29_v1;
wire                valid_24_to_29_v0,	valid_24_to_29_v1;
wire                ready_29_to_24_v0,	ready_29_to_24_v1;
wire    [`DW-1:0]   data_29_to_34_v0,	data_29_to_34_v1;
wire                valid_29_to_34_v0,	valid_29_to_34_v1;
wire                ready_34_to_29_v0,	ready_34_to_29_v1;
wire    [`DW-1:0]   data_34_to_39_v0,	data_34_to_39_v1;
wire                valid_34_to_39_v0,	valid_34_to_39_v1;
wire                ready_39_to_34_v0,	ready_39_to_34_v1;
wire    [`DW-1:0]   data_39_to_44_v0,	data_39_to_44_v1;
wire                valid_39_to_44_v0,	valid_39_to_44_v1;
wire                ready_44_to_39_v0,	ready_44_to_39_v1;
wire    [`DW-1:0]   data_44_to_49_v0,	data_44_to_49_v1;
wire                valid_44_to_49_v0,	valid_44_to_49_v1;
wire                ready_49_to_44_v0,	ready_49_to_44_v1;

/*Router 0,0*/    
cast_router #(
    .isUBM_list            (isUBM_list_0_0),
    .isFC_list             (isFC_list_0_0),
    .FCdn_list             (FCdn_list_0_0),
    .FCpl_list             (FCpl_list_0_0),
    .rt_file_list          (cast_rt_file_list_0_0)
)router_0_0(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_i_stab),
    .west_valid_i          (valid_i_stab),
    .west_ready_o          (ready_o_stab),
    .west_data_o           (),
    .west_valid_o          (),
    .west_ready_i          (1'b0),
    .east_data_i           (data_1_to_0),
    .east_valid_i          (valid_1_to_0),
    .east_ready_o          (ready_0_to_1),
    .east_data_o           (data_0_to_1),
    .east_valid_o          (valid_0_to_1),
    .east_ready_i          (ready_1_to_0),
    .vert0_data_i          (34'b0),
    .vert0_valid_i         (1'b0),
    .vert0_ready_o         (),
    .vert0_data_o          (data_0_to_5_v0),
    .vert0_valid_o         (valid_0_to_5_v0),
    .vert0_ready_i         (ready_5_to_0_v0),
    .vert1_data_i          (34'b0),
    .vert1_valid_i         (1'b0),
    .vert1_ready_o         (),
    .vert1_data_o          (data_0_to_5_v1),
    .vert1_valid_o         (valid_0_to_5_v1),
    .vert1_ready_i         (ready_5_to_0_v1),
    .local_data_i          (data_i[0][0]),
    .local_valid_i         (valid_i[0][0]),
    .local_ready_o         (ready_o[0][0]),
    .local_data_o          (data_o[0][0]),
    .local_valid_o         (valid_o[0][0]),
    .local_ready_i         (ready_i[0][0]),
    .credit_upd            (credit_upd)
);

/*Router 0,1*/    
cast_router #(
    .isUBM_list            (isUBM_list_0_1),
    .isFC_list             (isFC_list_0_1),
    .FCdn_list             (FCdn_list_0_1),
    .FCpl_list             (FCpl_list_0_1),
    .rt_file_list          (cast_rt_file_list_0_1)
)router_0_1(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (34'b0),
    .west_valid_i          (1'b0),
    .west_ready_o          (),
    .west_data_o           (),
    .west_valid_o          (),
    .west_ready_i          (1'b0),
    .east_data_i           (data_6_to_5),
    .east_valid_i          (valid_6_to_5),
    .east_ready_o          (ready_5_to_6),
    .east_data_o           (data_5_to_6),
    .east_valid_o          (valid_5_to_6),
    .east_ready_i          (ready_6_to_5),
    .vert0_data_i          (data_0_to_5_v0),
    .vert0_valid_i         (valid_0_to_5_v0),
    .vert0_ready_o         (ready_5_to_0_v0),
    .vert0_data_o          (data_5_to_10_v0),
    .vert0_valid_o         (valid_5_to_10_v0),
    .vert0_ready_i         (ready_10_to_5_v0),
    .vert1_data_i          (data_0_to_5_v1),
    .vert1_valid_i         (valid_0_to_5_v1),
    .vert1_ready_o         (ready_5_to_0_v1),
    .vert1_data_o          (data_5_to_10_v1),
    .vert1_valid_o         (valid_5_to_10_v1),
    .vert1_ready_i         (ready_10_to_5_v1),
    .local_data_i          (data_i[0][1]),
    .local_valid_i         (valid_i[0][1]),
    .local_ready_o         (ready_o[0][1]),
    .local_data_o          (data_o[0][1]),
    .local_valid_o         (valid_o[0][1]),
    .local_ready_i         (ready_i[0][1]),
    .credit_upd            (credit_upd)
);

/*Router 0,2*/    
cast_router #(
    .isUBM_list            (isUBM_list_0_2),
    .isFC_list             (isFC_list_0_2),
    .FCdn_list             (FCdn_list_0_2),
    .FCpl_list             (FCpl_list_0_2),
    .rt_file_list          (cast_rt_file_list_0_2)
)router_0_2(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (34'b0),
    .west_valid_i          (1'b0),
    .west_ready_o          (),
    .west_data_o           (),
    .west_valid_o          (),
    .west_ready_i          (1'b0),
    .east_data_i           (data_11_to_10),
    .east_valid_i          (valid_11_to_10),
    .east_ready_o          (ready_10_to_11),
    .east_data_o           (data_10_to_11),
    .east_valid_o          (valid_10_to_11),
    .east_ready_i          (ready_11_to_10),
    .vert0_data_i          (data_5_to_10_v0),
    .vert0_valid_i         (valid_5_to_10_v0),
    .vert0_ready_o         (ready_10_to_5_v0),
    .vert0_data_o          (data_10_to_15_v0),
    .vert0_valid_o         (valid_10_to_15_v0),
    .vert0_ready_i         (ready_15_to_10_v0),
    .vert1_data_i          (data_5_to_10_v1),
    .vert1_valid_i         (valid_5_to_10_v1),
    .vert1_ready_o         (ready_10_to_5_v1),
    .vert1_data_o          (data_10_to_15_v1),
    .vert1_valid_o         (valid_10_to_15_v1),
    .vert1_ready_i         (ready_15_to_10_v1),
    .local_data_i          (data_i[0][2]),
    .local_valid_i         (valid_i[0][2]),
    .local_ready_o         (ready_o[0][2]),
    .local_data_o          (data_o[0][2]),
    .local_valid_o         (valid_o[0][2]),
    .local_ready_i         (ready_i[0][2]),
    .credit_upd            (credit_upd)
);

/*Router 0,3*/    
cast_router #(
    .isUBM_list            (isUBM_list_0_3),
    .isFC_list             (isFC_list_0_3),
    .FCdn_list             (FCdn_list_0_3),
    .FCpl_list             (FCpl_list_0_3),
    .rt_file_list          (cast_rt_file_list_0_3)
)router_0_3(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (34'b0),
    .west_valid_i          (1'b0),
    .west_ready_o          (),
    .west_data_o           (),
    .west_valid_o          (),
    .west_ready_i          (1'b0),
    .east_data_i           (data_16_to_15),
    .east_valid_i          (valid_16_to_15),
    .east_ready_o          (ready_15_to_16),
    .east_data_o           (data_15_to_16),
    .east_valid_o          (valid_15_to_16),
    .east_ready_i          (ready_16_to_15),
    .vert0_data_i          (data_10_to_15_v0),
    .vert0_valid_i         (valid_10_to_15_v0),
    .vert0_ready_o         (ready_15_to_10_v0),
    .vert0_data_o          (data_15_to_20_v0),
    .vert0_valid_o         (valid_15_to_20_v0),
    .vert0_ready_i         (ready_20_to_15_v0),
    .vert1_data_i          (data_10_to_15_v1),
    .vert1_valid_i         (valid_10_to_15_v1),
    .vert1_ready_o         (ready_15_to_10_v1),
    .vert1_data_o          (data_15_to_20_v1),
    .vert1_valid_o         (valid_15_to_20_v1),
    .vert1_ready_i         (ready_20_to_15_v1),
    .local_data_i          (data_i[0][3]),
    .local_valid_i         (valid_i[0][3]),
    .local_ready_o         (ready_o[0][3]),
    .local_data_o          (data_o[0][3]),
    .local_valid_o         (valid_o[0][3]),
    .local_ready_i         (ready_i[0][3]),
    .credit_upd            (credit_upd)
);

/*Router 0,4*/    
cast_router #(
    .isUBM_list            (isUBM_list_0_4),
    .isFC_list             (isFC_list_0_4),
    .FCdn_list             (FCdn_list_0_4),
    .FCpl_list             (FCpl_list_0_4),
    .rt_file_list          (cast_rt_file_list_0_4)
)router_0_4(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (34'b0),
    .west_valid_i          (1'b0),
    .west_ready_o          (),
    .west_data_o           (),
    .west_valid_o          (),
    .west_ready_i          (1'b0),
    .east_data_i           (data_21_to_20),
    .east_valid_i          (valid_21_to_20),
    .east_ready_o          (ready_20_to_21),
    .east_data_o           (data_20_to_21),
    .east_valid_o          (valid_20_to_21),
    .east_ready_i          (ready_21_to_20),
    .vert0_data_i          (data_15_to_20_v0),
    .vert0_valid_i         (valid_15_to_20_v0),
    .vert0_ready_o         (ready_20_to_15_v0),
    .vert0_data_o          (data_20_to_25_v0),
    .vert0_valid_o         (valid_20_to_25_v0),
    .vert0_ready_i         (ready_25_to_20_v0),
    .vert1_data_i          (data_15_to_20_v1),
    .vert1_valid_i         (valid_15_to_20_v1),
    .vert1_ready_o         (ready_20_to_15_v1),
    .vert1_data_o          (data_20_to_25_v1),
    .vert1_valid_o         (valid_20_to_25_v1),
    .vert1_ready_i         (ready_25_to_20_v1),
    .local_data_i          (data_i[0][4]),
    .local_valid_i         (valid_i[0][4]),
    .local_ready_o         (ready_o[0][4]),
    .local_data_o          (data_o[0][4]),
    .local_valid_o         (valid_o[0][4]),
    .local_ready_i         (ready_i[0][4]),
    .credit_upd            (credit_upd)
);

/*Router 0,5*/    
cast_router #(
    .isUBM_list            (isUBM_list_0_5),
    .isFC_list             (isFC_list_0_5),
    .FCdn_list             (FCdn_list_0_5),
    .FCpl_list             (FCpl_list_0_5),
    .rt_file_list          (cast_rt_file_list_0_5)
)router_0_5(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (34'b0),
    .west_valid_i          (1'b0),
    .west_ready_o          (),
    .west_data_o           (),
    .west_valid_o          (),
    .west_ready_i          (1'b0),
    .east_data_i           (data_26_to_25),
    .east_valid_i          (valid_26_to_25),
    .east_ready_o          (ready_25_to_26),
    .east_data_o           (data_25_to_26),
    .east_valid_o          (valid_25_to_26),
    .east_ready_i          (ready_26_to_25),
    .vert0_data_i          (data_20_to_25_v0),
    .vert0_valid_i         (valid_20_to_25_v0),
    .vert0_ready_o         (ready_25_to_20_v0),
    .vert0_data_o          (data_25_to_30_v0),
    .vert0_valid_o         (valid_25_to_30_v0),
    .vert0_ready_i         (ready_30_to_25_v0),
    .vert1_data_i          (data_20_to_25_v1),
    .vert1_valid_i         (valid_20_to_25_v1),
    .vert1_ready_o         (ready_25_to_20_v1),
    .vert1_data_o          (data_25_to_30_v1),
    .vert1_valid_o         (valid_25_to_30_v1),
    .vert1_ready_i         (ready_30_to_25_v1),
    .local_data_i          (data_i[0][5]),
    .local_valid_i         (valid_i[0][5]),
    .local_ready_o         (ready_o[0][5]),
    .local_data_o          (data_o[0][5]),
    .local_valid_o         (valid_o[0][5]),
    .local_ready_i         (ready_i[0][5]),
    .credit_upd            (credit_upd)
);

/*Router 0,6*/    
cast_router #(
    .isUBM_list            (isUBM_list_0_6),
    .isFC_list             (isFC_list_0_6),
    .FCdn_list             (FCdn_list_0_6),
    .FCpl_list             (FCpl_list_0_6),
    .rt_file_list          (cast_rt_file_list_0_6)
)router_0_6(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (34'b0),
    .west_valid_i          (1'b0),
    .west_ready_o          (),
    .west_data_o           (),
    .west_valid_o          (),
    .west_ready_i          (1'b0),
    .east_data_i           (data_31_to_30),
    .east_valid_i          (valid_31_to_30),
    .east_ready_o          (ready_30_to_31),
    .east_data_o           (data_30_to_31),
    .east_valid_o          (valid_30_to_31),
    .east_ready_i          (ready_31_to_30),
    .vert0_data_i          (data_25_to_30_v0),
    .vert0_valid_i         (valid_25_to_30_v0),
    .vert0_ready_o         (ready_30_to_25_v0),
    .vert0_data_o          (data_30_to_35_v0),
    .vert0_valid_o         (valid_30_to_35_v0),
    .vert0_ready_i         (ready_35_to_30_v0),
    .vert1_data_i          (data_25_to_30_v1),
    .vert1_valid_i         (valid_25_to_30_v1),
    .vert1_ready_o         (ready_30_to_25_v1),
    .vert1_data_o          (data_30_to_35_v1),
    .vert1_valid_o         (valid_30_to_35_v1),
    .vert1_ready_i         (ready_35_to_30_v1),
    .local_data_i          (data_i[0][6]),
    .local_valid_i         (valid_i[0][6]),
    .local_ready_o         (ready_o[0][6]),
    .local_data_o          (data_o[0][6]),
    .local_valid_o         (valid_o[0][6]),
    .local_ready_i         (ready_i[0][6]),
    .credit_upd            (credit_upd)
);

/*Router 0,7*/    
cast_router #(
    .isUBM_list            (isUBM_list_0_7),
    .isFC_list             (isFC_list_0_7),
    .FCdn_list             (FCdn_list_0_7),
    .FCpl_list             (FCpl_list_0_7),
    .rt_file_list          (cast_rt_file_list_0_7)
)router_0_7(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (34'b0),
    .west_valid_i          (1'b0),
    .west_ready_o          (),
    .west_data_o           (),
    .west_valid_o          (),
    .west_ready_i          (1'b0),
    .east_data_i           (data_36_to_35),
    .east_valid_i          (valid_36_to_35),
    .east_ready_o          (ready_35_to_36),
    .east_data_o           (data_35_to_36),
    .east_valid_o          (valid_35_to_36),
    .east_ready_i          (ready_36_to_35),
    .vert0_data_i          (data_30_to_35_v0),
    .vert0_valid_i         (valid_30_to_35_v0),
    .vert0_ready_o         (ready_35_to_30_v0),
    .vert0_data_o          (data_35_to_40_v0),
    .vert0_valid_o         (valid_35_to_40_v0),
    .vert0_ready_i         (ready_40_to_35_v0),
    .vert1_data_i          (data_30_to_35_v1),
    .vert1_valid_i         (valid_30_to_35_v1),
    .vert1_ready_o         (ready_35_to_30_v1),
    .vert1_data_o          (data_35_to_40_v1),
    .vert1_valid_o         (valid_35_to_40_v1),
    .vert1_ready_i         (ready_40_to_35_v1),
    .local_data_i          (data_i[0][7]),
    .local_valid_i         (valid_i[0][7]),
    .local_ready_o         (ready_o[0][7]),
    .local_data_o          (data_o[0][7]),
    .local_valid_o         (valid_o[0][7]),
    .local_ready_i         (ready_i[0][7]),
    .credit_upd            (credit_upd)
);

/*Router 0,8*/    
cast_router #(
    .isUBM_list            (isUBM_list_0_8),
    .isFC_list             (isFC_list_0_8),
    .FCdn_list             (FCdn_list_0_8),
    .FCpl_list             (FCpl_list_0_8),
    .rt_file_list          (cast_rt_file_list_0_8)
)router_0_8(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (34'b0),
    .west_valid_i          (1'b0),
    .west_ready_o          (),
    .west_data_o           (),
    .west_valid_o          (),
    .west_ready_i          (1'b0),
    .east_data_i           (data_41_to_40),
    .east_valid_i          (valid_41_to_40),
    .east_ready_o          (ready_40_to_41),
    .east_data_o           (data_40_to_41),
    .east_valid_o          (valid_40_to_41),
    .east_ready_i          (ready_41_to_40),
    .vert0_data_i          (data_35_to_40_v0),
    .vert0_valid_i         (valid_35_to_40_v0),
    .vert0_ready_o         (ready_40_to_35_v0),
    .vert0_data_o          (data_40_to_45_v0),
    .vert0_valid_o         (valid_40_to_45_v0),
    .vert0_ready_i         (ready_45_to_40_v0),
    .vert1_data_i          (data_35_to_40_v1),
    .vert1_valid_i         (valid_35_to_40_v1),
    .vert1_ready_o         (ready_40_to_35_v1),
    .vert1_data_o          (data_40_to_45_v1),
    .vert1_valid_o         (valid_40_to_45_v1),
    .vert1_ready_i         (ready_45_to_40_v1),
    .local_data_i          (data_i[0][8]),
    .local_valid_i         (valid_i[0][8]),
    .local_ready_o         (ready_o[0][8]),
    .local_data_o          (data_o[0][8]),
    .local_valid_o         (valid_o[0][8]),
    .local_ready_i         (ready_i[0][8]),
    .credit_upd            (credit_upd)
);

/*Router 0,9*/    
cast_router #(
    .isUBM_list            (isUBM_list_0_9),
    .isFC_list             (isFC_list_0_9),
    .FCdn_list             (FCdn_list_0_9),
    .FCpl_list             (FCpl_list_0_9),
    .rt_file_list          (cast_rt_file_list_0_9)
)router_0_9(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (34'b0),
    .west_valid_i          (1'b0),
    .west_ready_o          (),
    .west_data_o           (),
    .west_valid_o          (),
    .west_ready_i          (1'b0),
    .east_data_i           (data_46_to_45),
    .east_valid_i          (valid_46_to_45),
    .east_ready_o          (ready_45_to_46),
    .east_data_o           (data_45_to_46),
    .east_valid_o          (valid_45_to_46),
    .east_ready_i          (ready_46_to_45),
    .vert0_data_i          (data_40_to_45_v0),
    .vert0_valid_i         (valid_40_to_45_v0),
    .vert0_ready_o         (ready_45_to_40_v0),
    .vert0_data_o          (),
    .vert0_valid_o         (),
    .vert0_ready_i         (1'b0),
    .vert1_data_i          (data_40_to_45_v1),
    .vert1_valid_i         (valid_40_to_45_v1),
    .vert1_ready_o         (ready_45_to_40_v1),
    .vert1_data_o          (),
    .vert1_valid_o         (),
    .vert1_ready_i         (1'b0),
    .local_data_i          (data_i[0][9]),
    .local_valid_i         (valid_i[0][9]),
    .local_ready_o         (ready_o[0][9]),
    .local_data_o          (data_o[0][9]),
    .local_valid_o         (valid_o[0][9]),
    .local_ready_i         (ready_i[0][9]),
    .credit_upd            (credit_upd)
);

/*Router 1,0*/    
cast_router #(
    .isUBM_list            (isUBM_list_1_0),
    .isFC_list             (isFC_list_1_0),
    .FCdn_list             (FCdn_list_1_0),
    .FCpl_list             (FCpl_list_1_0),
    .rt_file_list          (cast_rt_file_list_1_0)
)router_1_0(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_0_to_1),
    .west_valid_i          (valid_0_to_1),
    .west_ready_o          (ready_1_to_0),
    .west_data_o           (data_1_to_0),
    .west_valid_o          (valid_1_to_0),
    .west_ready_i          (ready_0_to_1),
    .east_data_i           (data_2_to_1),
    .east_valid_i          (valid_2_to_1),
    .east_ready_o          (ready_1_to_2),
    .east_data_o           (data_1_to_2),
    .east_valid_o          (valid_1_to_2),
    .east_ready_i          (ready_2_to_1),
    .vert0_data_i          (34'b0),
    .vert0_valid_i         (1'b0),
    .vert0_ready_o         (),
    .vert0_data_o          (data_1_to_6_v0),
    .vert0_valid_o         (valid_1_to_6_v0),
    .vert0_ready_i         (ready_6_to_1_v0),
    .vert1_data_i          (34'b0),
    .vert1_valid_i         (1'b0),
    .vert1_ready_o         (),
    .vert1_data_o          (data_1_to_6_v1),
    .vert1_valid_o         (valid_1_to_6_v1),
    .vert1_ready_i         (ready_6_to_1_v1),
    .local_data_i          (data_i[1][0]),
    .local_valid_i         (valid_i[1][0]),
    .local_ready_o         (ready_o[1][0]),
    .local_data_o          (data_o[1][0]),
    .local_valid_o         (valid_o[1][0]),
    .local_ready_i         (ready_i[1][0]),
    .credit_upd            (credit_upd)
);

/*Router 1,1*/    
cast_router #(
    .isUBM_list            (isUBM_list_1_1),
    .isFC_list             (isFC_list_1_1),
    .FCdn_list             (FCdn_list_1_1),
    .FCpl_list             (FCpl_list_1_1),
    .rt_file_list          (cast_rt_file_list_1_1)
)router_1_1(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_5_to_6),
    .west_valid_i          (valid_5_to_6),
    .west_ready_o          (ready_6_to_5),
    .west_data_o           (data_6_to_5),
    .west_valid_o          (valid_6_to_5),
    .west_ready_i          (ready_5_to_6),
    .east_data_i           (data_7_to_6),
    .east_valid_i          (valid_7_to_6),
    .east_ready_o          (ready_6_to_7),
    .east_data_o           (data_6_to_7),
    .east_valid_o          (valid_6_to_7),
    .east_ready_i          (ready_7_to_6),
    .vert0_data_i          (data_1_to_6_v0),
    .vert0_valid_i         (valid_1_to_6_v0),
    .vert0_ready_o         (ready_6_to_1_v0),
    .vert0_data_o          (data_6_to_11_v0),
    .vert0_valid_o         (valid_6_to_11_v0),
    .vert0_ready_i         (ready_11_to_6_v0),
    .vert1_data_i          (data_1_to_6_v1),
    .vert1_valid_i         (valid_1_to_6_v1),
    .vert1_ready_o         (ready_6_to_1_v1),
    .vert1_data_o          (data_6_to_11_v1),
    .vert1_valid_o         (valid_6_to_11_v1),
    .vert1_ready_i         (ready_11_to_6_v1),
    .local_data_i          (data_i[1][1]),
    .local_valid_i         (valid_i[1][1]),
    .local_ready_o         (ready_o[1][1]),
    .local_data_o          (data_o[1][1]),
    .local_valid_o         (valid_o[1][1]),
    .local_ready_i         (ready_i[1][1]),
    .credit_upd            (credit_upd)
);

/*Router 1,2*/    
cast_router #(
    .isUBM_list            (isUBM_list_1_2),
    .isFC_list             (isFC_list_1_2),
    .FCdn_list             (FCdn_list_1_2),
    .FCpl_list             (FCpl_list_1_2),
    .rt_file_list          (cast_rt_file_list_1_2)
)router_1_2(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_10_to_11),
    .west_valid_i          (valid_10_to_11),
    .west_ready_o          (ready_11_to_10),
    .west_data_o           (data_11_to_10),
    .west_valid_o          (valid_11_to_10),
    .west_ready_i          (ready_10_to_11),
    .east_data_i           (data_12_to_11),
    .east_valid_i          (valid_12_to_11),
    .east_ready_o          (ready_11_to_12),
    .east_data_o           (data_11_to_12),
    .east_valid_o          (valid_11_to_12),
    .east_ready_i          (ready_12_to_11),
    .vert0_data_i          (data_6_to_11_v0),
    .vert0_valid_i         (valid_6_to_11_v0),
    .vert0_ready_o         (ready_11_to_6_v0),
    .vert0_data_o          (data_11_to_16_v0),
    .vert0_valid_o         (valid_11_to_16_v0),
    .vert0_ready_i         (ready_16_to_11_v0),
    .vert1_data_i          (data_6_to_11_v1),
    .vert1_valid_i         (valid_6_to_11_v1),
    .vert1_ready_o         (ready_11_to_6_v1),
    .vert1_data_o          (data_11_to_16_v1),
    .vert1_valid_o         (valid_11_to_16_v1),
    .vert1_ready_i         (ready_16_to_11_v1),
    .local_data_i          (data_i[1][2]),
    .local_valid_i         (valid_i[1][2]),
    .local_ready_o         (ready_o[1][2]),
    .local_data_o          (data_o[1][2]),
    .local_valid_o         (valid_o[1][2]),
    .local_ready_i         (ready_i[1][2]),
    .credit_upd            (credit_upd)
);

/*Router 1,3*/    
cast_router #(
    .isUBM_list            (isUBM_list_1_3),
    .isFC_list             (isFC_list_1_3),
    .FCdn_list             (FCdn_list_1_3),
    .FCpl_list             (FCpl_list_1_3),
    .rt_file_list          (cast_rt_file_list_1_3)
)router_1_3(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_15_to_16),
    .west_valid_i          (valid_15_to_16),
    .west_ready_o          (ready_16_to_15),
    .west_data_o           (data_16_to_15),
    .west_valid_o          (valid_16_to_15),
    .west_ready_i          (ready_15_to_16),
    .east_data_i           (data_17_to_16),
    .east_valid_i          (valid_17_to_16),
    .east_ready_o          (ready_16_to_17),
    .east_data_o           (data_16_to_17),
    .east_valid_o          (valid_16_to_17),
    .east_ready_i          (ready_17_to_16),
    .vert0_data_i          (data_11_to_16_v0),
    .vert0_valid_i         (valid_11_to_16_v0),
    .vert0_ready_o         (ready_16_to_11_v0),
    .vert0_data_o          (data_16_to_21_v0),
    .vert0_valid_o         (valid_16_to_21_v0),
    .vert0_ready_i         (ready_21_to_16_v0),
    .vert1_data_i          (data_11_to_16_v1),
    .vert1_valid_i         (valid_11_to_16_v1),
    .vert1_ready_o         (ready_16_to_11_v1),
    .vert1_data_o          (data_16_to_21_v1),
    .vert1_valid_o         (valid_16_to_21_v1),
    .vert1_ready_i         (ready_21_to_16_v1),
    .local_data_i          (data_i[1][3]),
    .local_valid_i         (valid_i[1][3]),
    .local_ready_o         (ready_o[1][3]),
    .local_data_o          (data_o[1][3]),
    .local_valid_o         (valid_o[1][3]),
    .local_ready_i         (ready_i[1][3]),
    .credit_upd            (credit_upd)
);

/*Router 1,4*/    
cast_router #(
    .isUBM_list            (isUBM_list_1_4),
    .isFC_list             (isFC_list_1_4),
    .FCdn_list             (FCdn_list_1_4),
    .FCpl_list             (FCpl_list_1_4),
    .rt_file_list          (cast_rt_file_list_1_4)
)router_1_4(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_20_to_21),
    .west_valid_i          (valid_20_to_21),
    .west_ready_o          (ready_21_to_20),
    .west_data_o           (data_21_to_20),
    .west_valid_o          (valid_21_to_20),
    .west_ready_i          (ready_20_to_21),
    .east_data_i           (data_22_to_21),
    .east_valid_i          (valid_22_to_21),
    .east_ready_o          (ready_21_to_22),
    .east_data_o           (data_21_to_22),
    .east_valid_o          (valid_21_to_22),
    .east_ready_i          (ready_22_to_21),
    .vert0_data_i          (data_16_to_21_v0),
    .vert0_valid_i         (valid_16_to_21_v0),
    .vert0_ready_o         (ready_21_to_16_v0),
    .vert0_data_o          (data_21_to_26_v0),
    .vert0_valid_o         (valid_21_to_26_v0),
    .vert0_ready_i         (ready_26_to_21_v0),
    .vert1_data_i          (data_16_to_21_v1),
    .vert1_valid_i         (valid_16_to_21_v1),
    .vert1_ready_o         (ready_21_to_16_v1),
    .vert1_data_o          (data_21_to_26_v1),
    .vert1_valid_o         (valid_21_to_26_v1),
    .vert1_ready_i         (ready_26_to_21_v1),
    .local_data_i          (data_i[1][4]),
    .local_valid_i         (valid_i[1][4]),
    .local_ready_o         (ready_o[1][4]),
    .local_data_o          (data_o[1][4]),
    .local_valid_o         (valid_o[1][4]),
    .local_ready_i         (ready_i[1][4]),
    .credit_upd            (credit_upd)
);

/*Router 1,5*/    
cast_router #(
    .isUBM_list            (isUBM_list_1_5),
    .isFC_list             (isFC_list_1_5),
    .FCdn_list             (FCdn_list_1_5),
    .FCpl_list             (FCpl_list_1_5),
    .rt_file_list          (cast_rt_file_list_1_5)
)router_1_5(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_25_to_26),
    .west_valid_i          (valid_25_to_26),
    .west_ready_o          (ready_26_to_25),
    .west_data_o           (data_26_to_25),
    .west_valid_o          (valid_26_to_25),
    .west_ready_i          (ready_25_to_26),
    .east_data_i           (data_27_to_26),
    .east_valid_i          (valid_27_to_26),
    .east_ready_o          (ready_26_to_27),
    .east_data_o           (data_26_to_27),
    .east_valid_o          (valid_26_to_27),
    .east_ready_i          (ready_27_to_26),
    .vert0_data_i          (data_21_to_26_v0),
    .vert0_valid_i         (valid_21_to_26_v0),
    .vert0_ready_o         (ready_26_to_21_v0),
    .vert0_data_o          (data_26_to_31_v0),
    .vert0_valid_o         (valid_26_to_31_v0),
    .vert0_ready_i         (ready_31_to_26_v0),
    .vert1_data_i          (data_21_to_26_v1),
    .vert1_valid_i         (valid_21_to_26_v1),
    .vert1_ready_o         (ready_26_to_21_v1),
    .vert1_data_o          (data_26_to_31_v1),
    .vert1_valid_o         (valid_26_to_31_v1),
    .vert1_ready_i         (ready_31_to_26_v1),
    .local_data_i          (data_i[1][5]),
    .local_valid_i         (valid_i[1][5]),
    .local_ready_o         (ready_o[1][5]),
    .local_data_o          (data_o[1][5]),
    .local_valid_o         (valid_o[1][5]),
    .local_ready_i         (ready_i[1][5]),
    .credit_upd            (credit_upd)
);

/*Router 1,6*/    
cast_router #(
    .isUBM_list            (isUBM_list_1_6),
    .isFC_list             (isFC_list_1_6),
    .FCdn_list             (FCdn_list_1_6),
    .FCpl_list             (FCpl_list_1_6),
    .rt_file_list          (cast_rt_file_list_1_6)
)router_1_6(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_30_to_31),
    .west_valid_i          (valid_30_to_31),
    .west_ready_o          (ready_31_to_30),
    .west_data_o           (data_31_to_30),
    .west_valid_o          (valid_31_to_30),
    .west_ready_i          (ready_30_to_31),
    .east_data_i           (data_32_to_31),
    .east_valid_i          (valid_32_to_31),
    .east_ready_o          (ready_31_to_32),
    .east_data_o           (data_31_to_32),
    .east_valid_o          (valid_31_to_32),
    .east_ready_i          (ready_32_to_31),
    .vert0_data_i          (data_26_to_31_v0),
    .vert0_valid_i         (valid_26_to_31_v0),
    .vert0_ready_o         (ready_31_to_26_v0),
    .vert0_data_o          (data_31_to_36_v0),
    .vert0_valid_o         (valid_31_to_36_v0),
    .vert0_ready_i         (ready_36_to_31_v0),
    .vert1_data_i          (data_26_to_31_v1),
    .vert1_valid_i         (valid_26_to_31_v1),
    .vert1_ready_o         (ready_31_to_26_v1),
    .vert1_data_o          (data_31_to_36_v1),
    .vert1_valid_o         (valid_31_to_36_v1),
    .vert1_ready_i         (ready_36_to_31_v1),
    .local_data_i          (data_i[1][6]),
    .local_valid_i         (valid_i[1][6]),
    .local_ready_o         (ready_o[1][6]),
    .local_data_o          (data_o[1][6]),
    .local_valid_o         (valid_o[1][6]),
    .local_ready_i         (ready_i[1][6]),
    .credit_upd            (credit_upd)
);

/*Router 1,7*/    
cast_router #(
    .isUBM_list            (isUBM_list_1_7),
    .isFC_list             (isFC_list_1_7),
    .FCdn_list             (FCdn_list_1_7),
    .FCpl_list             (FCpl_list_1_7),
    .rt_file_list          (cast_rt_file_list_1_7)
)router_1_7(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_35_to_36),
    .west_valid_i          (valid_35_to_36),
    .west_ready_o          (ready_36_to_35),
    .west_data_o           (data_36_to_35),
    .west_valid_o          (valid_36_to_35),
    .west_ready_i          (ready_35_to_36),
    .east_data_i           (data_37_to_36),
    .east_valid_i          (valid_37_to_36),
    .east_ready_o          (ready_36_to_37),
    .east_data_o           (data_36_to_37),
    .east_valid_o          (valid_36_to_37),
    .east_ready_i          (ready_37_to_36),
    .vert0_data_i          (data_31_to_36_v0),
    .vert0_valid_i         (valid_31_to_36_v0),
    .vert0_ready_o         (ready_36_to_31_v0),
    .vert0_data_o          (data_36_to_41_v0),
    .vert0_valid_o         (valid_36_to_41_v0),
    .vert0_ready_i         (ready_41_to_36_v0),
    .vert1_data_i          (data_31_to_36_v1),
    .vert1_valid_i         (valid_31_to_36_v1),
    .vert1_ready_o         (ready_36_to_31_v1),
    .vert1_data_o          (data_36_to_41_v1),
    .vert1_valid_o         (valid_36_to_41_v1),
    .vert1_ready_i         (ready_41_to_36_v1),
    .local_data_i          (data_i[1][7]),
    .local_valid_i         (valid_i[1][7]),
    .local_ready_o         (ready_o[1][7]),
    .local_data_o          (data_o[1][7]),
    .local_valid_o         (valid_o[1][7]),
    .local_ready_i         (ready_i[1][7]),
    .credit_upd            (credit_upd)
);

/*Router 1,8*/    
cast_router #(
    .isUBM_list            (isUBM_list_1_8),
    .isFC_list             (isFC_list_1_8),
    .FCdn_list             (FCdn_list_1_8),
    .FCpl_list             (FCpl_list_1_8),
    .rt_file_list          (cast_rt_file_list_1_8)
)router_1_8(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_40_to_41),
    .west_valid_i          (valid_40_to_41),
    .west_ready_o          (ready_41_to_40),
    .west_data_o           (data_41_to_40),
    .west_valid_o          (valid_41_to_40),
    .west_ready_i          (ready_40_to_41),
    .east_data_i           (data_42_to_41),
    .east_valid_i          (valid_42_to_41),
    .east_ready_o          (ready_41_to_42),
    .east_data_o           (data_41_to_42),
    .east_valid_o          (valid_41_to_42),
    .east_ready_i          (ready_42_to_41),
    .vert0_data_i          (data_36_to_41_v0),
    .vert0_valid_i         (valid_36_to_41_v0),
    .vert0_ready_o         (ready_41_to_36_v0),
    .vert0_data_o          (data_41_to_46_v0),
    .vert0_valid_o         (valid_41_to_46_v0),
    .vert0_ready_i         (ready_46_to_41_v0),
    .vert1_data_i          (data_36_to_41_v1),
    .vert1_valid_i         (valid_36_to_41_v1),
    .vert1_ready_o         (ready_41_to_36_v1),
    .vert1_data_o          (data_41_to_46_v1),
    .vert1_valid_o         (valid_41_to_46_v1),
    .vert1_ready_i         (ready_46_to_41_v1),
    .local_data_i          (data_i[1][8]),
    .local_valid_i         (valid_i[1][8]),
    .local_ready_o         (ready_o[1][8]),
    .local_data_o          (data_o[1][8]),
    .local_valid_o         (valid_o[1][8]),
    .local_ready_i         (ready_i[1][8]),
    .credit_upd            (credit_upd)
);

/*Router 1,9*/    
cast_router #(
    .isUBM_list            (isUBM_list_1_9),
    .isFC_list             (isFC_list_1_9),
    .FCdn_list             (FCdn_list_1_9),
    .FCpl_list             (FCpl_list_1_9),
    .rt_file_list          (cast_rt_file_list_1_9)
)router_1_9(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_45_to_46),
    .west_valid_i          (valid_45_to_46),
    .west_ready_o          (ready_46_to_45),
    .west_data_o           (data_46_to_45),
    .west_valid_o          (valid_46_to_45),
    .west_ready_i          (ready_45_to_46),
    .east_data_i           (data_47_to_46),
    .east_valid_i          (valid_47_to_46),
    .east_ready_o          (ready_46_to_47),
    .east_data_o           (data_46_to_47),
    .east_valid_o          (valid_46_to_47),
    .east_ready_i          (ready_47_to_46),
    .vert0_data_i          (data_41_to_46_v0),
    .vert0_valid_i         (valid_41_to_46_v0),
    .vert0_ready_o         (ready_46_to_41_v0),
    .vert0_data_o          (),
    .vert0_valid_o         (),
    .vert0_ready_i         (1'b0),
    .vert1_data_i          (data_41_to_46_v1),
    .vert1_valid_i         (valid_41_to_46_v1),
    .vert1_ready_o         (ready_46_to_41_v1),
    .vert1_data_o          (),
    .vert1_valid_o         (),
    .vert1_ready_i         (1'b0),
    .local_data_i          (data_i[1][9]),
    .local_valid_i         (valid_i[1][9]),
    .local_ready_o         (ready_o[1][9]),
    .local_data_o          (data_o[1][9]),
    .local_valid_o         (valid_o[1][9]),
    .local_ready_i         (ready_i[1][9]),
    .credit_upd            (credit_upd)
);

/*Router 2,0*/    
cast_router #(
    .isUBM_list            (isUBM_list_2_0),
    .isFC_list             (isFC_list_2_0),
    .FCdn_list             (FCdn_list_2_0),
    .FCpl_list             (FCpl_list_2_0),
    .rt_file_list          (cast_rt_file_list_2_0)
)router_2_0(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_1_to_2),
    .west_valid_i          (valid_1_to_2),
    .west_ready_o          (ready_2_to_1),
    .west_data_o           (data_2_to_1),
    .west_valid_o          (valid_2_to_1),
    .west_ready_i          (ready_1_to_2),
    .east_data_i           (data_3_to_2),
    .east_valid_i          (valid_3_to_2),
    .east_ready_o          (ready_2_to_3),
    .east_data_o           (data_2_to_3),
    .east_valid_o          (valid_2_to_3),
    .east_ready_i          (ready_3_to_2),
    .vert0_data_i          (34'b0),
    .vert0_valid_i         (1'b0),
    .vert0_ready_o         (),
    .vert0_data_o          (data_2_to_7_v0),
    .vert0_valid_o         (valid_2_to_7_v0),
    .vert0_ready_i         (ready_7_to_2_v0),
    .vert1_data_i          (34'b0),
    .vert1_valid_i         (1'b0),
    .vert1_ready_o         (),
    .vert1_data_o          (data_2_to_7_v1),
    .vert1_valid_o         (valid_2_to_7_v1),
    .vert1_ready_i         (ready_7_to_2_v1),
    .local_data_i          (data_i[2][0]),
    .local_valid_i         (valid_i[2][0]),
    .local_ready_o         (ready_o[2][0]),
    .local_data_o          (data_o[2][0]),
    .local_valid_o         (valid_o[2][0]),
    .local_ready_i         (ready_i[2][0]),
    .credit_upd            (credit_upd)
);

/*Router 2,1*/    
cast_router #(
    .isUBM_list            (isUBM_list_2_1),
    .isFC_list             (isFC_list_2_1),
    .FCdn_list             (FCdn_list_2_1),
    .FCpl_list             (FCpl_list_2_1),
    .rt_file_list          (cast_rt_file_list_2_1)
)router_2_1(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_6_to_7),
    .west_valid_i          (valid_6_to_7),
    .west_ready_o          (ready_7_to_6),
    .west_data_o           (data_7_to_6),
    .west_valid_o          (valid_7_to_6),
    .west_ready_i          (ready_6_to_7),
    .east_data_i           (data_8_to_7),
    .east_valid_i          (valid_8_to_7),
    .east_ready_o          (ready_7_to_8),
    .east_data_o           (data_7_to_8),
    .east_valid_o          (valid_7_to_8),
    .east_ready_i          (ready_8_to_7),
    .vert0_data_i          (data_2_to_7_v0),
    .vert0_valid_i         (valid_2_to_7_v0),
    .vert0_ready_o         (ready_7_to_2_v0),
    .vert0_data_o          (data_7_to_12_v0),
    .vert0_valid_o         (valid_7_to_12_v0),
    .vert0_ready_i         (ready_12_to_7_v0),
    .vert1_data_i          (data_2_to_7_v1),
    .vert1_valid_i         (valid_2_to_7_v1),
    .vert1_ready_o         (ready_7_to_2_v1),
    .vert1_data_o          (data_7_to_12_v1),
    .vert1_valid_o         (valid_7_to_12_v1),
    .vert1_ready_i         (ready_12_to_7_v1),
    .local_data_i          (data_i[2][1]),
    .local_valid_i         (valid_i[2][1]),
    .local_ready_o         (ready_o[2][1]),
    .local_data_o          (data_o[2][1]),
    .local_valid_o         (valid_o[2][1]),
    .local_ready_i         (ready_i[2][1]),
    .credit_upd            (credit_upd)
);

/*Router 2,2*/    
cast_router #(
    .isUBM_list            (isUBM_list_2_2),
    .isFC_list             (isFC_list_2_2),
    .FCdn_list             (FCdn_list_2_2),
    .FCpl_list             (FCpl_list_2_2),
    .rt_file_list          (cast_rt_file_list_2_2)
)router_2_2(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_11_to_12),
    .west_valid_i          (valid_11_to_12),
    .west_ready_o          (ready_12_to_11),
    .west_data_o           (data_12_to_11),
    .west_valid_o          (valid_12_to_11),
    .west_ready_i          (ready_11_to_12),
    .east_data_i           (data_13_to_12),
    .east_valid_i          (valid_13_to_12),
    .east_ready_o          (ready_12_to_13),
    .east_data_o           (data_12_to_13),
    .east_valid_o          (valid_12_to_13),
    .east_ready_i          (ready_13_to_12),
    .vert0_data_i          (data_7_to_12_v0),
    .vert0_valid_i         (valid_7_to_12_v0),
    .vert0_ready_o         (ready_12_to_7_v0),
    .vert0_data_o          (data_12_to_17_v0),
    .vert0_valid_o         (valid_12_to_17_v0),
    .vert0_ready_i         (ready_17_to_12_v0),
    .vert1_data_i          (data_7_to_12_v1),
    .vert1_valid_i         (valid_7_to_12_v1),
    .vert1_ready_o         (ready_12_to_7_v1),
    .vert1_data_o          (data_12_to_17_v1),
    .vert1_valid_o         (valid_12_to_17_v1),
    .vert1_ready_i         (ready_17_to_12_v1),
    .local_data_i          (data_i[2][2]),
    .local_valid_i         (valid_i[2][2]),
    .local_ready_o         (ready_o[2][2]),
    .local_data_o          (data_o[2][2]),
    .local_valid_o         (valid_o[2][2]),
    .local_ready_i         (ready_i[2][2]),
    .credit_upd            (credit_upd)
);

/*Router 2,3*/    
cast_router #(
    .isUBM_list            (isUBM_list_2_3),
    .isFC_list             (isFC_list_2_3),
    .FCdn_list             (FCdn_list_2_3),
    .FCpl_list             (FCpl_list_2_3),
    .rt_file_list          (cast_rt_file_list_2_3)
)router_2_3(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_16_to_17),
    .west_valid_i          (valid_16_to_17),
    .west_ready_o          (ready_17_to_16),
    .west_data_o           (data_17_to_16),
    .west_valid_o          (valid_17_to_16),
    .west_ready_i          (ready_16_to_17),
    .east_data_i           (data_18_to_17),
    .east_valid_i          (valid_18_to_17),
    .east_ready_o          (ready_17_to_18),
    .east_data_o           (data_17_to_18),
    .east_valid_o          (valid_17_to_18),
    .east_ready_i          (ready_18_to_17),
    .vert0_data_i          (data_12_to_17_v0),
    .vert0_valid_i         (valid_12_to_17_v0),
    .vert0_ready_o         (ready_17_to_12_v0),
    .vert0_data_o          (data_17_to_22_v0),
    .vert0_valid_o         (valid_17_to_22_v0),
    .vert0_ready_i         (ready_22_to_17_v0),
    .vert1_data_i          (data_12_to_17_v1),
    .vert1_valid_i         (valid_12_to_17_v1),
    .vert1_ready_o         (ready_17_to_12_v1),
    .vert1_data_o          (data_17_to_22_v1),
    .vert1_valid_o         (valid_17_to_22_v1),
    .vert1_ready_i         (ready_22_to_17_v1),
    .local_data_i          (data_i[2][3]),
    .local_valid_i         (valid_i[2][3]),
    .local_ready_o         (ready_o[2][3]),
    .local_data_o          (data_o[2][3]),
    .local_valid_o         (valid_o[2][3]),
    .local_ready_i         (ready_i[2][3]),
    .credit_upd            (credit_upd)
);

/*Router 2,4*/    
cast_router #(
    .isUBM_list            (isUBM_list_2_4),
    .isFC_list             (isFC_list_2_4),
    .FCdn_list             (FCdn_list_2_4),
    .FCpl_list             (FCpl_list_2_4),
    .rt_file_list          (cast_rt_file_list_2_4)
)router_2_4(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_21_to_22),
    .west_valid_i          (valid_21_to_22),
    .west_ready_o          (ready_22_to_21),
    .west_data_o           (data_22_to_21),
    .west_valid_o          (valid_22_to_21),
    .west_ready_i          (ready_21_to_22),
    .east_data_i           (data_23_to_22),
    .east_valid_i          (valid_23_to_22),
    .east_ready_o          (ready_22_to_23),
    .east_data_o           (data_22_to_23),
    .east_valid_o          (valid_22_to_23),
    .east_ready_i          (ready_23_to_22),
    .vert0_data_i          (data_17_to_22_v0),
    .vert0_valid_i         (valid_17_to_22_v0),
    .vert0_ready_o         (ready_22_to_17_v0),
    .vert0_data_o          (data_22_to_27_v0),
    .vert0_valid_o         (valid_22_to_27_v0),
    .vert0_ready_i         (ready_27_to_22_v0),
    .vert1_data_i          (data_17_to_22_v1),
    .vert1_valid_i         (valid_17_to_22_v1),
    .vert1_ready_o         (ready_22_to_17_v1),
    .vert1_data_o          (data_22_to_27_v1),
    .vert1_valid_o         (valid_22_to_27_v1),
    .vert1_ready_i         (ready_27_to_22_v1),
    .local_data_i          (data_i[2][4]),
    .local_valid_i         (valid_i[2][4]),
    .local_ready_o         (ready_o[2][4]),
    .local_data_o          (data_o[2][4]),
    .local_valid_o         (valid_o[2][4]),
    .local_ready_i         (ready_i[2][4]),
    .credit_upd            (credit_upd)
);

/*Router 2,5*/    
cast_router #(
    .isUBM_list            (isUBM_list_2_5),
    .isFC_list             (isFC_list_2_5),
    .FCdn_list             (FCdn_list_2_5),
    .FCpl_list             (FCpl_list_2_5),
    .rt_file_list          (cast_rt_file_list_2_5)
)router_2_5(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_26_to_27),
    .west_valid_i          (valid_26_to_27),
    .west_ready_o          (ready_27_to_26),
    .west_data_o           (data_27_to_26),
    .west_valid_o          (valid_27_to_26),
    .west_ready_i          (ready_26_to_27),
    .east_data_i           (data_28_to_27),
    .east_valid_i          (valid_28_to_27),
    .east_ready_o          (ready_27_to_28),
    .east_data_o           (data_27_to_28),
    .east_valid_o          (valid_27_to_28),
    .east_ready_i          (ready_28_to_27),
    .vert0_data_i          (data_22_to_27_v0),
    .vert0_valid_i         (valid_22_to_27_v0),
    .vert0_ready_o         (ready_27_to_22_v0),
    .vert0_data_o          (data_27_to_32_v0),
    .vert0_valid_o         (valid_27_to_32_v0),
    .vert0_ready_i         (ready_32_to_27_v0),
    .vert1_data_i          (data_22_to_27_v1),
    .vert1_valid_i         (valid_22_to_27_v1),
    .vert1_ready_o         (ready_27_to_22_v1),
    .vert1_data_o          (data_27_to_32_v1),
    .vert1_valid_o         (valid_27_to_32_v1),
    .vert1_ready_i         (ready_32_to_27_v1),
    .local_data_i          (data_i[2][5]),
    .local_valid_i         (valid_i[2][5]),
    .local_ready_o         (ready_o[2][5]),
    .local_data_o          (data_o[2][5]),
    .local_valid_o         (valid_o[2][5]),
    .local_ready_i         (ready_i[2][5]),
    .credit_upd            (credit_upd)
);

/*Router 2,6*/    
cast_router #(
    .isUBM_list            (isUBM_list_2_6),
    .isFC_list             (isFC_list_2_6),
    .FCdn_list             (FCdn_list_2_6),
    .FCpl_list             (FCpl_list_2_6),
    .rt_file_list          (cast_rt_file_list_2_6)
)router_2_6(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_31_to_32),
    .west_valid_i          (valid_31_to_32),
    .west_ready_o          (ready_32_to_31),
    .west_data_o           (data_32_to_31),
    .west_valid_o          (valid_32_to_31),
    .west_ready_i          (ready_31_to_32),
    .east_data_i           (data_33_to_32),
    .east_valid_i          (valid_33_to_32),
    .east_ready_o          (ready_32_to_33),
    .east_data_o           (data_32_to_33),
    .east_valid_o          (valid_32_to_33),
    .east_ready_i          (ready_33_to_32),
    .vert0_data_i          (data_27_to_32_v0),
    .vert0_valid_i         (valid_27_to_32_v0),
    .vert0_ready_o         (ready_32_to_27_v0),
    .vert0_data_o          (data_32_to_37_v0),
    .vert0_valid_o         (valid_32_to_37_v0),
    .vert0_ready_i         (ready_37_to_32_v0),
    .vert1_data_i          (data_27_to_32_v1),
    .vert1_valid_i         (valid_27_to_32_v1),
    .vert1_ready_o         (ready_32_to_27_v1),
    .vert1_data_o          (data_32_to_37_v1),
    .vert1_valid_o         (valid_32_to_37_v1),
    .vert1_ready_i         (ready_37_to_32_v1),
    .local_data_i          (data_i[2][6]),
    .local_valid_i         (valid_i[2][6]),
    .local_ready_o         (ready_o[2][6]),
    .local_data_o          (data_o[2][6]),
    .local_valid_o         (valid_o[2][6]),
    .local_ready_i         (ready_i[2][6]),
    .credit_upd            (credit_upd)
);

/*Router 2,7*/    
cast_router #(
    .isUBM_list            (isUBM_list_2_7),
    .isFC_list             (isFC_list_2_7),
    .FCdn_list             (FCdn_list_2_7),
    .FCpl_list             (FCpl_list_2_7),
    .rt_file_list          (cast_rt_file_list_2_7)
)router_2_7(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_36_to_37),
    .west_valid_i          (valid_36_to_37),
    .west_ready_o          (ready_37_to_36),
    .west_data_o           (data_37_to_36),
    .west_valid_o          (valid_37_to_36),
    .west_ready_i          (ready_36_to_37),
    .east_data_i           (data_38_to_37),
    .east_valid_i          (valid_38_to_37),
    .east_ready_o          (ready_37_to_38),
    .east_data_o           (data_37_to_38),
    .east_valid_o          (valid_37_to_38),
    .east_ready_i          (ready_38_to_37),
    .vert0_data_i          (data_32_to_37_v0),
    .vert0_valid_i         (valid_32_to_37_v0),
    .vert0_ready_o         (ready_37_to_32_v0),
    .vert0_data_o          (data_37_to_42_v0),
    .vert0_valid_o         (valid_37_to_42_v0),
    .vert0_ready_i         (ready_42_to_37_v0),
    .vert1_data_i          (data_32_to_37_v1),
    .vert1_valid_i         (valid_32_to_37_v1),
    .vert1_ready_o         (ready_37_to_32_v1),
    .vert1_data_o          (data_37_to_42_v1),
    .vert1_valid_o         (valid_37_to_42_v1),
    .vert1_ready_i         (ready_42_to_37_v1),
    .local_data_i          (data_i[2][7]),
    .local_valid_i         (valid_i[2][7]),
    .local_ready_o         (ready_o[2][7]),
    .local_data_o          (data_o[2][7]),
    .local_valid_o         (valid_o[2][7]),
    .local_ready_i         (ready_i[2][7]),
    .credit_upd            (credit_upd)
);

/*Router 2,8*/    
cast_router #(
    .isUBM_list            (isUBM_list_2_8),
    .isFC_list             (isFC_list_2_8),
    .FCdn_list             (FCdn_list_2_8),
    .FCpl_list             (FCpl_list_2_8),
    .rt_file_list          (cast_rt_file_list_2_8)
)router_2_8(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_41_to_42),
    .west_valid_i          (valid_41_to_42),
    .west_ready_o          (ready_42_to_41),
    .west_data_o           (data_42_to_41),
    .west_valid_o          (valid_42_to_41),
    .west_ready_i          (ready_41_to_42),
    .east_data_i           (data_43_to_42),
    .east_valid_i          (valid_43_to_42),
    .east_ready_o          (ready_42_to_43),
    .east_data_o           (data_42_to_43),
    .east_valid_o          (valid_42_to_43),
    .east_ready_i          (ready_43_to_42),
    .vert0_data_i          (data_37_to_42_v0),
    .vert0_valid_i         (valid_37_to_42_v0),
    .vert0_ready_o         (ready_42_to_37_v0),
    .vert0_data_o          (data_42_to_47_v0),
    .vert0_valid_o         (valid_42_to_47_v0),
    .vert0_ready_i         (ready_47_to_42_v0),
    .vert1_data_i          (data_37_to_42_v1),
    .vert1_valid_i         (valid_37_to_42_v1),
    .vert1_ready_o         (ready_42_to_37_v1),
    .vert1_data_o          (data_42_to_47_v1),
    .vert1_valid_o         (valid_42_to_47_v1),
    .vert1_ready_i         (ready_47_to_42_v1),
    .local_data_i          (data_i[2][8]),
    .local_valid_i         (valid_i[2][8]),
    .local_ready_o         (ready_o[2][8]),
    .local_data_o          (data_o[2][8]),
    .local_valid_o         (valid_o[2][8]),
    .local_ready_i         (ready_i[2][8]),
    .credit_upd            (credit_upd)
);

/*Router 2,9*/    
cast_router #(
    .isUBM_list            (isUBM_list_2_9),
    .isFC_list             (isFC_list_2_9),
    .FCdn_list             (FCdn_list_2_9),
    .FCpl_list             (FCpl_list_2_9),
    .rt_file_list          (cast_rt_file_list_2_9)
)router_2_9(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_46_to_47),
    .west_valid_i          (valid_46_to_47),
    .west_ready_o          (ready_47_to_46),
    .west_data_o           (data_47_to_46),
    .west_valid_o          (valid_47_to_46),
    .west_ready_i          (ready_46_to_47),
    .east_data_i           (data_48_to_47),
    .east_valid_i          (valid_48_to_47),
    .east_ready_o          (ready_47_to_48),
    .east_data_o           (data_47_to_48),
    .east_valid_o          (valid_47_to_48),
    .east_ready_i          (ready_48_to_47),
    .vert0_data_i          (data_42_to_47_v0),
    .vert0_valid_i         (valid_42_to_47_v0),
    .vert0_ready_o         (ready_47_to_42_v0),
    .vert0_data_o          (),
    .vert0_valid_o         (),
    .vert0_ready_i         (1'b0),
    .vert1_data_i          (data_42_to_47_v1),
    .vert1_valid_i         (valid_42_to_47_v1),
    .vert1_ready_o         (ready_47_to_42_v1),
    .vert1_data_o          (),
    .vert1_valid_o         (),
    .vert1_ready_i         (1'b0),
    .local_data_i          (data_i[2][9]),
    .local_valid_i         (valid_i[2][9]),
    .local_ready_o         (ready_o[2][9]),
    .local_data_o          (data_o[2][9]),
    .local_valid_o         (valid_o[2][9]),
    .local_ready_i         (ready_i[2][9]),
    .credit_upd            (credit_upd)
);

/*Router 3,0*/    
cast_router #(
    .isUBM_list            (isUBM_list_3_0),
    .isFC_list             (isFC_list_3_0),
    .FCdn_list             (FCdn_list_3_0),
    .FCpl_list             (FCpl_list_3_0),
    .rt_file_list          (cast_rt_file_list_3_0)
)router_3_0(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_2_to_3),
    .west_valid_i          (valid_2_to_3),
    .west_ready_o          (ready_3_to_2),
    .west_data_o           (data_3_to_2),
    .west_valid_o          (valid_3_to_2),
    .west_ready_i          (ready_2_to_3),
    .east_data_i           (data_4_to_3),
    .east_valid_i          (valid_4_to_3),
    .east_ready_o          (ready_3_to_4),
    .east_data_o           (data_3_to_4),
    .east_valid_o          (valid_3_to_4),
    .east_ready_i          (ready_4_to_3),
    .vert0_data_i          (34'b0),
    .vert0_valid_i         (1'b0),
    .vert0_ready_o         (),
    .vert0_data_o          (data_3_to_8_v0),
    .vert0_valid_o         (valid_3_to_8_v0),
    .vert0_ready_i         (ready_8_to_3_v0),
    .vert1_data_i          (34'b0),
    .vert1_valid_i         (1'b0),
    .vert1_ready_o         (),
    .vert1_data_o          (data_3_to_8_v1),
    .vert1_valid_o         (valid_3_to_8_v1),
    .vert1_ready_i         (ready_8_to_3_v1),
    .local_data_i          (data_i[3][0]),
    .local_valid_i         (valid_i[3][0]),
    .local_ready_o         (ready_o[3][0]),
    .local_data_o          (data_o[3][0]),
    .local_valid_o         (valid_o[3][0]),
    .local_ready_i         (ready_i[3][0]),
    .credit_upd            (credit_upd)
);

/*Router 3,1*/    
cast_router #(
    .isUBM_list            (isUBM_list_3_1),
    .isFC_list             (isFC_list_3_1),
    .FCdn_list             (FCdn_list_3_1),
    .FCpl_list             (FCpl_list_3_1),
    .rt_file_list          (cast_rt_file_list_3_1)
)router_3_1(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_7_to_8),
    .west_valid_i          (valid_7_to_8),
    .west_ready_o          (ready_8_to_7),
    .west_data_o           (data_8_to_7),
    .west_valid_o          (valid_8_to_7),
    .west_ready_i          (ready_7_to_8),
    .east_data_i           (data_9_to_8),
    .east_valid_i          (valid_9_to_8),
    .east_ready_o          (ready_8_to_9),
    .east_data_o           (data_8_to_9),
    .east_valid_o          (valid_8_to_9),
    .east_ready_i          (ready_9_to_8),
    .vert0_data_i          (data_3_to_8_v0),
    .vert0_valid_i         (valid_3_to_8_v0),
    .vert0_ready_o         (ready_8_to_3_v0),
    .vert0_data_o          (data_8_to_13_v0),
    .vert0_valid_o         (valid_8_to_13_v0),
    .vert0_ready_i         (ready_13_to_8_v0),
    .vert1_data_i          (data_3_to_8_v1),
    .vert1_valid_i         (valid_3_to_8_v1),
    .vert1_ready_o         (ready_8_to_3_v1),
    .vert1_data_o          (data_8_to_13_v1),
    .vert1_valid_o         (valid_8_to_13_v1),
    .vert1_ready_i         (ready_13_to_8_v1),
    .local_data_i          (data_i[3][1]),
    .local_valid_i         (valid_i[3][1]),
    .local_ready_o         (ready_o[3][1]),
    .local_data_o          (data_o[3][1]),
    .local_valid_o         (valid_o[3][1]),
    .local_ready_i         (ready_i[3][1]),
    .credit_upd            (credit_upd)
);

/*Router 3,2*/    
cast_router #(
    .isUBM_list            (isUBM_list_3_2),
    .isFC_list             (isFC_list_3_2),
    .FCdn_list             (FCdn_list_3_2),
    .FCpl_list             (FCpl_list_3_2),
    .rt_file_list          (cast_rt_file_list_3_2)
)router_3_2(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_12_to_13),
    .west_valid_i          (valid_12_to_13),
    .west_ready_o          (ready_13_to_12),
    .west_data_o           (data_13_to_12),
    .west_valid_o          (valid_13_to_12),
    .west_ready_i          (ready_12_to_13),
    .east_data_i           (data_14_to_13),
    .east_valid_i          (valid_14_to_13),
    .east_ready_o          (ready_13_to_14),
    .east_data_o           (data_13_to_14),
    .east_valid_o          (valid_13_to_14),
    .east_ready_i          (ready_14_to_13),
    .vert0_data_i          (data_8_to_13_v0),
    .vert0_valid_i         (valid_8_to_13_v0),
    .vert0_ready_o         (ready_13_to_8_v0),
    .vert0_data_o          (data_13_to_18_v0),
    .vert0_valid_o         (valid_13_to_18_v0),
    .vert0_ready_i         (ready_18_to_13_v0),
    .vert1_data_i          (data_8_to_13_v1),
    .vert1_valid_i         (valid_8_to_13_v1),
    .vert1_ready_o         (ready_13_to_8_v1),
    .vert1_data_o          (data_13_to_18_v1),
    .vert1_valid_o         (valid_13_to_18_v1),
    .vert1_ready_i         (ready_18_to_13_v1),
    .local_data_i          (data_i[3][2]),
    .local_valid_i         (valid_i[3][2]),
    .local_ready_o         (ready_o[3][2]),
    .local_data_o          (data_o[3][2]),
    .local_valid_o         (valid_o[3][2]),
    .local_ready_i         (ready_i[3][2]),
    .credit_upd            (credit_upd)
);

/*Router 3,3*/    
cast_router #(
    .isUBM_list            (isUBM_list_3_3),
    .isFC_list             (isFC_list_3_3),
    .FCdn_list             (FCdn_list_3_3),
    .FCpl_list             (FCpl_list_3_3),
    .rt_file_list          (cast_rt_file_list_3_3)
)router_3_3(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_17_to_18),
    .west_valid_i          (valid_17_to_18),
    .west_ready_o          (ready_18_to_17),
    .west_data_o           (data_18_to_17),
    .west_valid_o          (valid_18_to_17),
    .west_ready_i          (ready_17_to_18),
    .east_data_i           (data_19_to_18),
    .east_valid_i          (valid_19_to_18),
    .east_ready_o          (ready_18_to_19),
    .east_data_o           (data_18_to_19),
    .east_valid_o          (valid_18_to_19),
    .east_ready_i          (ready_19_to_18),
    .vert0_data_i          (data_13_to_18_v0),
    .vert0_valid_i         (valid_13_to_18_v0),
    .vert0_ready_o         (ready_18_to_13_v0),
    .vert0_data_o          (data_18_to_23_v0),
    .vert0_valid_o         (valid_18_to_23_v0),
    .vert0_ready_i         (ready_23_to_18_v0),
    .vert1_data_i          (data_13_to_18_v1),
    .vert1_valid_i         (valid_13_to_18_v1),
    .vert1_ready_o         (ready_18_to_13_v1),
    .vert1_data_o          (data_18_to_23_v1),
    .vert1_valid_o         (valid_18_to_23_v1),
    .vert1_ready_i         (ready_23_to_18_v1),
    .local_data_i          (data_i[3][3]),
    .local_valid_i         (valid_i[3][3]),
    .local_ready_o         (ready_o[3][3]),
    .local_data_o          (data_o[3][3]),
    .local_valid_o         (valid_o[3][3]),
    .local_ready_i         (ready_i[3][3]),
    .credit_upd            (credit_upd)
);

/*Router 3,4*/    
cast_router #(
    .isUBM_list            (isUBM_list_3_4),
    .isFC_list             (isFC_list_3_4),
    .FCdn_list             (FCdn_list_3_4),
    .FCpl_list             (FCpl_list_3_4),
    .rt_file_list          (cast_rt_file_list_3_4)
)router_3_4(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_22_to_23),
    .west_valid_i          (valid_22_to_23),
    .west_ready_o          (ready_23_to_22),
    .west_data_o           (data_23_to_22),
    .west_valid_o          (valid_23_to_22),
    .west_ready_i          (ready_22_to_23),
    .east_data_i           (data_24_to_23),
    .east_valid_i          (valid_24_to_23),
    .east_ready_o          (ready_23_to_24),
    .east_data_o           (data_23_to_24),
    .east_valid_o          (valid_23_to_24),
    .east_ready_i          (ready_24_to_23),
    .vert0_data_i          (data_18_to_23_v0),
    .vert0_valid_i         (valid_18_to_23_v0),
    .vert0_ready_o         (ready_23_to_18_v0),
    .vert0_data_o          (data_23_to_28_v0),
    .vert0_valid_o         (valid_23_to_28_v0),
    .vert0_ready_i         (ready_28_to_23_v0),
    .vert1_data_i          (data_18_to_23_v1),
    .vert1_valid_i         (valid_18_to_23_v1),
    .vert1_ready_o         (ready_23_to_18_v1),
    .vert1_data_o          (data_23_to_28_v1),
    .vert1_valid_o         (valid_23_to_28_v1),
    .vert1_ready_i         (ready_28_to_23_v1),
    .local_data_i          (data_i[3][4]),
    .local_valid_i         (valid_i[3][4]),
    .local_ready_o         (ready_o[3][4]),
    .local_data_o          (data_o[3][4]),
    .local_valid_o         (valid_o[3][4]),
    .local_ready_i         (ready_i[3][4]),
    .credit_upd            (credit_upd)
);

/*Router 3,5*/    
cast_router #(
    .isUBM_list            (isUBM_list_3_5),
    .isFC_list             (isFC_list_3_5),
    .FCdn_list             (FCdn_list_3_5),
    .FCpl_list             (FCpl_list_3_5),
    .rt_file_list          (cast_rt_file_list_3_5)
)router_3_5(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_27_to_28),
    .west_valid_i          (valid_27_to_28),
    .west_ready_o          (ready_28_to_27),
    .west_data_o           (data_28_to_27),
    .west_valid_o          (valid_28_to_27),
    .west_ready_i          (ready_27_to_28),
    .east_data_i           (data_29_to_28),
    .east_valid_i          (valid_29_to_28),
    .east_ready_o          (ready_28_to_29),
    .east_data_o           (data_28_to_29),
    .east_valid_o          (valid_28_to_29),
    .east_ready_i          (ready_29_to_28),
    .vert0_data_i          (data_23_to_28_v0),
    .vert0_valid_i         (valid_23_to_28_v0),
    .vert0_ready_o         (ready_28_to_23_v0),
    .vert0_data_o          (data_28_to_33_v0),
    .vert0_valid_o         (valid_28_to_33_v0),
    .vert0_ready_i         (ready_33_to_28_v0),
    .vert1_data_i          (data_23_to_28_v1),
    .vert1_valid_i         (valid_23_to_28_v1),
    .vert1_ready_o         (ready_28_to_23_v1),
    .vert1_data_o          (data_28_to_33_v1),
    .vert1_valid_o         (valid_28_to_33_v1),
    .vert1_ready_i         (ready_33_to_28_v1),
    .local_data_i          (data_i[3][5]),
    .local_valid_i         (valid_i[3][5]),
    .local_ready_o         (ready_o[3][5]),
    .local_data_o          (data_o[3][5]),
    .local_valid_o         (valid_o[3][5]),
    .local_ready_i         (ready_i[3][5]),
    .credit_upd            (credit_upd)
);

/*Router 3,6*/    
cast_router #(
    .isUBM_list            (isUBM_list_3_6),
    .isFC_list             (isFC_list_3_6),
    .FCdn_list             (FCdn_list_3_6),
    .FCpl_list             (FCpl_list_3_6),
    .rt_file_list          (cast_rt_file_list_3_6)
)router_3_6(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_32_to_33),
    .west_valid_i          (valid_32_to_33),
    .west_ready_o          (ready_33_to_32),
    .west_data_o           (data_33_to_32),
    .west_valid_o          (valid_33_to_32),
    .west_ready_i          (ready_32_to_33),
    .east_data_i           (data_34_to_33),
    .east_valid_i          (valid_34_to_33),
    .east_ready_o          (ready_33_to_34),
    .east_data_o           (data_33_to_34),
    .east_valid_o          (valid_33_to_34),
    .east_ready_i          (ready_34_to_33),
    .vert0_data_i          (data_28_to_33_v0),
    .vert0_valid_i         (valid_28_to_33_v0),
    .vert0_ready_o         (ready_33_to_28_v0),
    .vert0_data_o          (data_33_to_38_v0),
    .vert0_valid_o         (valid_33_to_38_v0),
    .vert0_ready_i         (ready_38_to_33_v0),
    .vert1_data_i          (data_28_to_33_v1),
    .vert1_valid_i         (valid_28_to_33_v1),
    .vert1_ready_o         (ready_33_to_28_v1),
    .vert1_data_o          (data_33_to_38_v1),
    .vert1_valid_o         (valid_33_to_38_v1),
    .vert1_ready_i         (ready_38_to_33_v1),
    .local_data_i          (data_i[3][6]),
    .local_valid_i         (valid_i[3][6]),
    .local_ready_o         (ready_o[3][6]),
    .local_data_o          (data_o[3][6]),
    .local_valid_o         (valid_o[3][6]),
    .local_ready_i         (ready_i[3][6]),
    .credit_upd            (credit_upd)
);

/*Router 3,7*/    
cast_router #(
    .isUBM_list            (isUBM_list_3_7),
    .isFC_list             (isFC_list_3_7),
    .FCdn_list             (FCdn_list_3_7),
    .FCpl_list             (FCpl_list_3_7),
    .rt_file_list          (cast_rt_file_list_3_7)
)router_3_7(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_37_to_38),
    .west_valid_i          (valid_37_to_38),
    .west_ready_o          (ready_38_to_37),
    .west_data_o           (data_38_to_37),
    .west_valid_o          (valid_38_to_37),
    .west_ready_i          (ready_37_to_38),
    .east_data_i           (data_39_to_38),
    .east_valid_i          (valid_39_to_38),
    .east_ready_o          (ready_38_to_39),
    .east_data_o           (data_38_to_39),
    .east_valid_o          (valid_38_to_39),
    .east_ready_i          (ready_39_to_38),
    .vert0_data_i          (data_33_to_38_v0),
    .vert0_valid_i         (valid_33_to_38_v0),
    .vert0_ready_o         (ready_38_to_33_v0),
    .vert0_data_o          (data_38_to_43_v0),
    .vert0_valid_o         (valid_38_to_43_v0),
    .vert0_ready_i         (ready_43_to_38_v0),
    .vert1_data_i          (data_33_to_38_v1),
    .vert1_valid_i         (valid_33_to_38_v1),
    .vert1_ready_o         (ready_38_to_33_v1),
    .vert1_data_o          (data_38_to_43_v1),
    .vert1_valid_o         (valid_38_to_43_v1),
    .vert1_ready_i         (ready_43_to_38_v1),
    .local_data_i          (data_i[3][7]),
    .local_valid_i         (valid_i[3][7]),
    .local_ready_o         (ready_o[3][7]),
    .local_data_o          (data_o[3][7]),
    .local_valid_o         (valid_o[3][7]),
    .local_ready_i         (ready_i[3][7]),
    .credit_upd            (credit_upd)
);

/*Router 3,8*/    
cast_router #(
    .isUBM_list            (isUBM_list_3_8),
    .isFC_list             (isFC_list_3_8),
    .FCdn_list             (FCdn_list_3_8),
    .FCpl_list             (FCpl_list_3_8),
    .rt_file_list          (cast_rt_file_list_3_8)
)router_3_8(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_42_to_43),
    .west_valid_i          (valid_42_to_43),
    .west_ready_o          (ready_43_to_42),
    .west_data_o           (data_43_to_42),
    .west_valid_o          (valid_43_to_42),
    .west_ready_i          (ready_42_to_43),
    .east_data_i           (data_44_to_43),
    .east_valid_i          (valid_44_to_43),
    .east_ready_o          (ready_43_to_44),
    .east_data_o           (data_o_flee00),
    .east_valid_o          (valid_o_flee0),
    .east_ready_i          (ready_i_flee0),
    .vert0_data_i          (data_38_to_43_v0),
    .vert0_valid_i         (valid_38_to_43_v0),
    .vert0_ready_o         (ready_43_to_38_v0),
    .vert0_data_o          (data_43_to_48_v0),
    .vert0_valid_o         (valid_43_to_48_v0),
    .vert0_ready_i         (ready_48_to_43_v0),
    .vert1_data_i          (data_38_to_43_v1),
    .vert1_valid_i         (valid_38_to_43_v1),
    .vert1_ready_o         (ready_43_to_38_v1),
    .vert1_data_o          (data_43_to_48_v1),
    .vert1_valid_o         (valid_43_to_48_v1),
    .vert1_ready_i         (ready_48_to_43_v1),
    .local_data_i          (data_i[3][8]),
    .local_valid_i         (valid_i[3][8]),
    .local_ready_o         (ready_o[3][8]),
    .local_data_o          (data_o[3][8]),
    .local_valid_o         (valid_o[3][8]),
    .local_ready_i         (ready_i[3][8]),
    .credit_upd            (credit_upd)
);

/*Router 3,9*/    
cast_router #(
    .isUBM_list            (isUBM_list_3_9),
    .isFC_list             (isFC_list_3_9),
    .FCdn_list             (FCdn_list_3_9),
    .FCpl_list             (FCpl_list_3_9),
    .rt_file_list          (cast_rt_file_list_3_9)
)router_3_9(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_47_to_48),
    .west_valid_i          (valid_47_to_48),
    .west_ready_o          (ready_48_to_47),
    .west_data_o           (data_o_flee1),
    .west_valid_o          (valid_o_flee1),
    .west_ready_i          (ready_i_flee1),
    .east_data_i           (data_49_to_48),
    .east_valid_i          (valid_49_to_48),
    .east_ready_o          (ready_48_to_49),
    .east_data_o           (data_48_to_49),
    .east_valid_o          (valid_48_to_49),
    .east_ready_i          (ready_49_to_48),
    .vert0_data_i          (data_43_to_48_v0),
    .vert0_valid_i         (valid_43_to_48_v0),
    .vert0_ready_o         (ready_48_to_43_v0),
    .vert0_data_o          (),
    .vert0_valid_o         (),
    .vert0_ready_i         (1'b0),
    .vert1_data_i          (data_43_to_48_v1),
    .vert1_valid_i         (valid_43_to_48_v1),
    .vert1_ready_o         (ready_48_to_43_v1),
    .vert1_data_o          (),
    .vert1_valid_o         (),
    .vert1_ready_i         (1'b0),
    .local_data_i          (data_i[3][9]),
    .local_valid_i         (valid_i[3][9]),
    .local_ready_o         (ready_o[3][9]),
    .local_data_o          (data_o[3][9]),
    .local_valid_o         (valid_o[3][9]),
    .local_ready_i         (ready_i[3][9]),
    .credit_upd            (credit_upd)
);

/*Router 4,0*/    
cast_router #(
    .isUBM_list            (isUBM_list_4_0),
    .isFC_list             (isFC_list_4_0),
    .FCdn_list             (FCdn_list_4_0),
    .FCpl_list             (FCpl_list_4_0),
    .rt_file_list          (cast_rt_file_list_4_0)
)router_4_0(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_3_to_4),
    .west_valid_i          (valid_3_to_4),
    .west_ready_o          (ready_4_to_3),
    .west_data_o           (data_4_to_3),
    .west_valid_o          (valid_4_to_3),
    .west_ready_i          (ready_3_to_4),
    .east_data_i           (34'b0),
    .east_valid_i          (1'b0),
    .east_ready_o          (),
    .east_data_o           (),
    .east_valid_o          (),
    .east_ready_i          (1'b0),
    .vert0_data_i          (34'b0),
    .vert0_valid_i         (1'b0),
    .vert0_ready_o         (),
    .vert0_data_o          (data_4_to_9_v0),
    .vert0_valid_o         (valid_4_to_9_v0),
    .vert0_ready_i         (ready_9_to_4_v0),
    .vert1_data_i          (34'b0),
    .vert1_valid_i         (1'b0),
    .vert1_ready_o         (),
    .vert1_data_o          (data_4_to_9_v1),
    .vert1_valid_o         (valid_4_to_9_v1),
    .vert1_ready_i         (ready_9_to_4_v1),
    .local_data_i          (data_i[4][0]),
    .local_valid_i         (valid_i[4][0]),
    .local_ready_o         (ready_o[4][0]),
    .local_data_o          (data_o[4][0]),
    .local_valid_o         (valid_o[4][0]),
    .local_ready_i         (ready_i[4][0]),
    .credit_upd            (credit_upd)
);

/*Router 4,1*/    
cast_router #(
    .isUBM_list            (isUBM_list_4_1),
    .isFC_list             (isFC_list_4_1),
    .FCdn_list             (FCdn_list_4_1),
    .FCpl_list             (FCpl_list_4_1),
    .rt_file_list          (cast_rt_file_list_4_1)
)router_4_1(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_8_to_9),
    .west_valid_i          (valid_8_to_9),
    .west_ready_o          (ready_9_to_8),
    .west_data_o           (data_9_to_8),
    .west_valid_o          (valid_9_to_8),
    .west_ready_i          (ready_8_to_9),
    .east_data_i           (34'b0),
    .east_valid_i          (1'b0),
    .east_ready_o          (),
    .east_data_o           (),
    .east_valid_o          (),
    .east_ready_i          (1'b0),
    .vert0_data_i          (data_4_to_9_v0),
    .vert0_valid_i         (valid_4_to_9_v0),
    .vert0_ready_o         (ready_9_to_4_v0),
    .vert0_data_o          (data_9_to_14_v0),
    .vert0_valid_o         (valid_9_to_14_v0),
    .vert0_ready_i         (ready_14_to_9_v0),
    .vert1_data_i          (data_4_to_9_v1),
    .vert1_valid_i         (valid_4_to_9_v1),
    .vert1_ready_o         (ready_9_to_4_v1),
    .vert1_data_o          (data_9_to_14_v1),
    .vert1_valid_o         (valid_9_to_14_v1),
    .vert1_ready_i         (ready_14_to_9_v1),
    .local_data_i          (data_i[4][1]),
    .local_valid_i         (valid_i[4][1]),
    .local_ready_o         (ready_o[4][1]),
    .local_data_o          (data_o[4][1]),
    .local_valid_o         (valid_o[4][1]),
    .local_ready_i         (ready_i[4][1]),
    .credit_upd            (credit_upd)
);

/*Router 4,2*/    
cast_router #(
    .isUBM_list            (isUBM_list_4_2),
    .isFC_list             (isFC_list_4_2),
    .FCdn_list             (FCdn_list_4_2),
    .FCpl_list             (FCpl_list_4_2),
    .rt_file_list          (cast_rt_file_list_4_2)
)router_4_2(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_13_to_14),
    .west_valid_i          (valid_13_to_14),
    .west_ready_o          (ready_14_to_13),
    .west_data_o           (data_14_to_13),
    .west_valid_o          (valid_14_to_13),
    .west_ready_i          (ready_13_to_14),
    .east_data_i           (34'b0),
    .east_valid_i          (1'b0),
    .east_ready_o          (),
    .east_data_o           (),
    .east_valid_o          (),
    .east_ready_i          (1'b0),
    .vert0_data_i          (data_9_to_14_v0),
    .vert0_valid_i         (valid_9_to_14_v0),
    .vert0_ready_o         (ready_14_to_9_v0),
    .vert0_data_o          (data_14_to_19_v0),
    .vert0_valid_o         (valid_14_to_19_v0),
    .vert0_ready_i         (ready_19_to_14_v0),
    .vert1_data_i          (data_9_to_14_v1),
    .vert1_valid_i         (valid_9_to_14_v1),
    .vert1_ready_o         (ready_14_to_9_v1),
    .vert1_data_o          (data_14_to_19_v1),
    .vert1_valid_o         (valid_14_to_19_v1),
    .vert1_ready_i         (ready_19_to_14_v1),
    .local_data_i          (data_i[4][2]),
    .local_valid_i         (valid_i[4][2]),
    .local_ready_o         (ready_o[4][2]),
    .local_data_o          (data_o[4][2]),
    .local_valid_o         (valid_o[4][2]),
    .local_ready_i         (ready_i[4][2]),
    .credit_upd            (credit_upd)
);

/*Router 4,3*/    
cast_router #(
    .isUBM_list            (isUBM_list_4_3),
    .isFC_list             (isFC_list_4_3),
    .FCdn_list             (FCdn_list_4_3),
    .FCpl_list             (FCpl_list_4_3),
    .rt_file_list          (cast_rt_file_list_4_3)
)router_4_3(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_18_to_19),
    .west_valid_i          (valid_18_to_19),
    .west_ready_o          (ready_19_to_18),
    .west_data_o           (data_19_to_18),
    .west_valid_o          (valid_19_to_18),
    .west_ready_i          (ready_18_to_19),
    .east_data_i           (34'b0),
    .east_valid_i          (1'b0),
    .east_ready_o          (),
    .east_data_o           (),
    .east_valid_o          (),
    .east_ready_i          (1'b0),
    .vert0_data_i          (data_14_to_19_v0),
    .vert0_valid_i         (valid_14_to_19_v0),
    .vert0_ready_o         (ready_19_to_14_v0),
    .vert0_data_o          (data_19_to_24_v0),
    .vert0_valid_o         (valid_19_to_24_v0),
    .vert0_ready_i         (ready_24_to_19_v0),
    .vert1_data_i          (data_14_to_19_v1),
    .vert1_valid_i         (valid_14_to_19_v1),
    .vert1_ready_o         (ready_19_to_14_v1),
    .vert1_data_o          (data_19_to_24_v1),
    .vert1_valid_o         (valid_19_to_24_v1),
    .vert1_ready_i         (ready_24_to_19_v1),
    .local_data_i          (data_i[4][3]),
    .local_valid_i         (valid_i[4][3]),
    .local_ready_o         (ready_o[4][3]),
    .local_data_o          (data_o[4][3]),
    .local_valid_o         (valid_o[4][3]),
    .local_ready_i         (ready_i[4][3]),
    .credit_upd            (credit_upd)
);

/*Router 4,4*/    
cast_router #(
    .isUBM_list            (isUBM_list_4_4),
    .isFC_list             (isFC_list_4_4),
    .FCdn_list             (FCdn_list_4_4),
    .FCpl_list             (FCpl_list_4_4),
    .rt_file_list          (cast_rt_file_list_4_4)
)router_4_4(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_23_to_24),
    .west_valid_i          (valid_23_to_24),
    .west_ready_o          (ready_24_to_23),
    .west_data_o           (data_24_to_23),
    .west_valid_o          (valid_24_to_23),
    .west_ready_i          (ready_23_to_24),
    .east_data_i           (34'b0),
    .east_valid_i          (1'b0),
    .east_ready_o          (),
    .east_data_o           (),
    .east_valid_o          (),
    .east_ready_i          (1'b0),
    .vert0_data_i          (data_19_to_24_v0),
    .vert0_valid_i         (valid_19_to_24_v0),
    .vert0_ready_o         (ready_24_to_19_v0),
    .vert0_data_o          (data_24_to_29_v0),
    .vert0_valid_o         (valid_24_to_29_v0),
    .vert0_ready_i         (ready_29_to_24_v0),
    .vert1_data_i          (data_19_to_24_v1),
    .vert1_valid_i         (valid_19_to_24_v1),
    .vert1_ready_o         (ready_24_to_19_v1),
    .vert1_data_o          (data_24_to_29_v1),
    .vert1_valid_o         (valid_24_to_29_v1),
    .vert1_ready_i         (ready_29_to_24_v1),
    .local_data_i          (data_i[4][4]),
    .local_valid_i         (valid_i[4][4]),
    .local_ready_o         (ready_o[4][4]),
    .local_data_o          (data_o[4][4]),
    .local_valid_o         (valid_o[4][4]),
    .local_ready_i         (ready_i[4][4]),
    .credit_upd            (credit_upd)
);

/*Router 4,5*/    
cast_router #(
    .isUBM_list            (isUBM_list_4_5),
    .isFC_list             (isFC_list_4_5),
    .FCdn_list             (FCdn_list_4_5),
    .FCpl_list             (FCpl_list_4_5),
    .rt_file_list          (cast_rt_file_list_4_5)
)router_4_5(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_28_to_29),
    .west_valid_i          (valid_28_to_29),
    .west_ready_o          (ready_29_to_28),
    .west_data_o           (data_29_to_28),
    .west_valid_o          (valid_29_to_28),
    .west_ready_i          (ready_28_to_29),
    .east_data_i           (34'b0),
    .east_valid_i          (1'b0),
    .east_ready_o          (),
    .east_data_o           (),
    .east_valid_o          (),
    .east_ready_i          (1'b0),
    .vert0_data_i          (data_24_to_29_v0),
    .vert0_valid_i         (valid_24_to_29_v0),
    .vert0_ready_o         (ready_29_to_24_v0),
    .vert0_data_o          (data_29_to_34_v0),
    .vert0_valid_o         (valid_29_to_34_v0),
    .vert0_ready_i         (ready_34_to_29_v0),
    .vert1_data_i          (data_24_to_29_v1),
    .vert1_valid_i         (valid_24_to_29_v1),
    .vert1_ready_o         (ready_29_to_24_v1),
    .vert1_data_o          (data_29_to_34_v1),
    .vert1_valid_o         (valid_29_to_34_v1),
    .vert1_ready_i         (ready_34_to_29_v1),
    .local_data_i          (data_i[4][5]),
    .local_valid_i         (valid_i[4][5]),
    .local_ready_o         (ready_o[4][5]),
    .local_data_o          (data_o[4][5]),
    .local_valid_o         (valid_o[4][5]),
    .local_ready_i         (ready_i[4][5]),
    .credit_upd            (credit_upd)
);

/*Router 4,6*/    
cast_router #(
    .isUBM_list            (isUBM_list_4_6),
    .isFC_list             (isFC_list_4_6),
    .FCdn_list             (FCdn_list_4_6),
    .FCpl_list             (FCpl_list_4_6),
    .rt_file_list          (cast_rt_file_list_4_6)
)router_4_6(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_33_to_34),
    .west_valid_i          (valid_33_to_34),
    .west_ready_o          (ready_34_to_33),
    .west_data_o           (data_34_to_33),
    .west_valid_o          (valid_34_to_33),
    .west_ready_i          (ready_33_to_34),
    .east_data_i           (34'b0),
    .east_valid_i          (1'b0),
    .east_ready_o          (),
    .east_data_o           (),
    .east_valid_o          (),
    .east_ready_i          (1'b0),
    .vert0_data_i          (data_29_to_34_v0),
    .vert0_valid_i         (valid_29_to_34_v0),
    .vert0_ready_o         (ready_34_to_29_v0),
    .vert0_data_o          (data_34_to_39_v0),
    .vert0_valid_o         (valid_34_to_39_v0),
    .vert0_ready_i         (ready_39_to_34_v0),
    .vert1_data_i          (data_29_to_34_v1),
    .vert1_valid_i         (valid_29_to_34_v1),
    .vert1_ready_o         (ready_34_to_29_v1),
    .vert1_data_o          (data_34_to_39_v1),
    .vert1_valid_o         (valid_34_to_39_v1),
    .vert1_ready_i         (ready_39_to_34_v1),
    .local_data_i          (data_i[4][6]),
    .local_valid_i         (valid_i[4][6]),
    .local_ready_o         (ready_o[4][6]),
    .local_data_o          (data_o[4][6]),
    .local_valid_o         (valid_o[4][6]),
    .local_ready_i         (ready_i[4][6]),
    .credit_upd            (credit_upd)
);

/*Router 4,7*/    
cast_router #(
    .isUBM_list            (isUBM_list_4_7),
    .isFC_list             (isFC_list_4_7),
    .FCdn_list             (FCdn_list_4_7),
    .FCpl_list             (FCpl_list_4_7),
    .rt_file_list          (cast_rt_file_list_4_7)
)router_4_7(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_38_to_39),
    .west_valid_i          (valid_38_to_39),
    .west_ready_o          (ready_39_to_38),
    .west_data_o           (data_39_to_38),
    .west_valid_o          (valid_39_to_38),
    .west_ready_i          (ready_38_to_39),
    .east_data_i           (34'b0),
    .east_valid_i          (1'b0),
    .east_ready_o          (),
    .east_data_o           (),
    .east_valid_o          (),
    .east_ready_i          (1'b0),
    .vert0_data_i          (data_34_to_39_v0),
    .vert0_valid_i         (valid_34_to_39_v0),
    .vert0_ready_o         (ready_39_to_34_v0),
    .vert0_data_o          (data_39_to_44_v0),
    .vert0_valid_o         (valid_39_to_44_v0),
    .vert0_ready_i         (ready_44_to_39_v0),
    .vert1_data_i          (data_34_to_39_v1),
    .vert1_valid_i         (valid_34_to_39_v1),
    .vert1_ready_o         (ready_39_to_34_v1),
    .vert1_data_o          (data_39_to_44_v1),
    .vert1_valid_o         (valid_39_to_44_v1),
    .vert1_ready_i         (ready_44_to_39_v1),
    .local_data_i          (data_i[4][7]),
    .local_valid_i         (valid_i[4][7]),
    .local_ready_o         (ready_o[4][7]),
    .local_data_o          (data_o[4][7]),
    .local_valid_o         (valid_o[4][7]),
    .local_ready_i         (ready_i[4][7]),
    .credit_upd            (credit_upd)
);

/*Router 4,8*/    
cast_router #(
    .isUBM_list            (isUBM_list_4_8),
    .isFC_list             (isFC_list_4_8),
    .FCdn_list             (FCdn_list_4_8),
    .FCpl_list             (FCpl_list_4_8),
    .rt_file_list          (cast_rt_file_list_4_8)
)router_4_8(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_43_to_44),
    .west_valid_i          (valid_43_to_44),
    .west_ready_o          (ready_44_to_43),
    .west_data_o           (data_44_to_43),
    .west_valid_o          (valid_44_to_43),
    .west_ready_i          (ready_43_to_44),
    .east_data_i           (34'b0),
    .east_valid_i          (1'b0),
    .east_ready_o          (),
    .east_data_o           (),
    .east_valid_o          (),
    .east_ready_i          (1'b0),
    .vert0_data_i          (data_39_to_44_v0),
    .vert0_valid_i         (valid_39_to_44_v0),
    .vert0_ready_o         (ready_44_to_39_v0),
    .vert0_data_o          (data_44_to_49_v0),
    .vert0_valid_o         (valid_44_to_49_v0),
    .vert0_ready_i         (ready_49_to_44_v0),
    .vert1_data_i          (data_39_to_44_v1),
    .vert1_valid_i         (valid_39_to_44_v1),
    .vert1_ready_o         (ready_44_to_39_v1),
    .vert1_data_o          (data_44_to_49_v1),
    .vert1_valid_o         (valid_44_to_49_v1),
    .vert1_ready_i         (ready_49_to_44_v1),
    .local_data_i          (data_i[4][8]),
    .local_valid_i         (valid_i[4][8]),
    .local_ready_o         (ready_o[4][8]),
    .local_data_o          (data_o[4][8]),
    .local_valid_o         (valid_o[4][8]),
    .local_ready_i         (ready_i[4][8]),
    .credit_upd            (credit_upd)
);

/*Router 4,9*/    
cast_router #(
    .isUBM_list            (isUBM_list_4_9),
    .isFC_list             (isFC_list_4_9),
    .FCdn_list             (FCdn_list_4_9),
    .FCpl_list             (FCpl_list_4_9),
    .rt_file_list          (cast_rt_file_list_4_9)
)router_4_9(
    .clk                   (clk),
    .rstn                  (rstn),
    .west_data_i           (data_48_to_49),
    .west_valid_i          (valid_48_to_49),
    .west_ready_o          (ready_49_to_48),
    .west_data_o           (data_49_to_48),
    .west_valid_o          (valid_49_to_48),
    .west_ready_i          (ready_48_to_49),
    .east_data_i           (34'b0),
    .east_valid_i          (1'b0),
    .east_ready_o          (),
    .east_data_o           (),
    .east_valid_o          (),
    .east_ready_i          (1'b0),
    .vert0_data_i          (data_44_to_49_v0),
    .vert0_valid_i         (valid_44_to_49_v0),
    .vert0_ready_o         (ready_49_to_44_v0),
    .vert0_data_o          (),
    .vert0_valid_o         (),
    .vert0_ready_i         (1'b0),
    .vert1_data_i          (data_44_to_49_v1),
    .vert1_valid_i         (valid_44_to_49_v1),
    .vert1_ready_o         (ready_49_to_44_v1),
    .vert1_data_o          (),
    .vert1_valid_o         (),
    .vert1_ready_i         (1'b0),
    .local_data_i          (data_i[4][9]),
    .local_valid_i         (valid_i[4][9]),
    .local_ready_o         (ready_o[4][9]),
    .local_data_o          (data_o[4][9]),
    .local_valid_o         (valid_o[4][9]),
    .local_ready_i         (ready_i[4][9]),
    .credit_upd            (credit_upd)
);

endmodule
