
`ifndef __GATHER_NETWORK_CONFIG_SVH_
`define __GATHER_NETWORK_CONFIG_SVH_
    
localparam string gather_rt_file_list_0_0[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_0_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_0_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_0_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_0_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_0_4"};

localparam string gather_rt_file_list_0_1[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_1_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_1_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_1_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_1_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_1_4"};

localparam string gather_rt_file_list_0_2[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_2_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_2_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_2_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_2_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_2_4"};

localparam string gather_rt_file_list_0_3[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_3_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_3_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_3_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_3_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_3_4"};

localparam string gather_rt_file_list_0_4[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_4_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_4_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_4_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_4_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_4_4"};

localparam string gather_rt_file_list_0_5[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_5_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_5_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_5_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_5_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_5_4"};

localparam string gather_rt_file_list_0_6[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_6_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_6_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_6_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_6_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_6_4"};

localparam string gather_rt_file_list_0_7[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_7_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_7_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_7_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_7_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_7_4"};

localparam string gather_rt_file_list_0_8[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_8_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_8_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_8_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_8_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_8_4"};

localparam string gather_rt_file_list_0_9[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_9_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_9_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_9_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_9_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_9_4"};

localparam string gather_rt_file_list_0_10[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_10_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_10_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_10_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_10_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_10_4"};

localparam string gather_rt_file_list_0_11[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_11_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_11_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_11_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_11_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_11_4"};

localparam string gather_rt_file_list_0_12[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_12_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_12_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_12_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_12_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_12_4"};

localparam string gather_rt_file_list_0_13[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_13_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_13_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_13_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_13_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_13_4"};

localparam string gather_rt_file_list_0_14[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_14_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_14_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_14_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_14_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_14_4"};

localparam string gather_rt_file_list_0_15[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_15_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_15_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_15_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_15_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_15_4"};

localparam string gather_rt_file_list_0_16[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_16_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_16_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_16_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_16_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_16_4"};

localparam string gather_rt_file_list_0_17[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_17_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_17_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_17_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_17_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_17_4"};

localparam string gather_rt_file_list_0_18[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_18_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_18_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_18_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_18_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_18_4"};

localparam string gather_rt_file_list_0_19[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_19_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_19_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_19_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_19_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_19_4"};

localparam string gather_rt_file_list_0_20[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_20_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_20_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_20_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_20_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_20_4"};

localparam string gather_rt_file_list_0_21[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_21_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_21_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_21_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_21_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_21_4"};

localparam string gather_rt_file_list_0_22[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_22_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_22_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_22_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_22_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_22_4"};

localparam string gather_rt_file_list_0_23[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_23_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_23_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_23_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_23_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_23_4"};

localparam string gather_rt_file_list_0_24[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_24_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_24_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_24_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_24_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_0_24_4"};

localparam string gather_rt_file_list_1_0[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_0_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_0_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_0_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_0_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_0_4"};

localparam string gather_rt_file_list_1_1[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_1_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_1_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_1_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_1_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_1_4"};

localparam string gather_rt_file_list_1_2[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_2_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_2_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_2_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_2_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_2_4"};

localparam string gather_rt_file_list_1_3[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_3_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_3_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_3_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_3_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_3_4"};

localparam string gather_rt_file_list_1_4[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_4_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_4_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_4_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_4_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_4_4"};

localparam string gather_rt_file_list_1_5[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_5_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_5_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_5_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_5_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_5_4"};

localparam string gather_rt_file_list_1_6[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_6_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_6_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_6_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_6_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_6_4"};

localparam string gather_rt_file_list_1_7[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_7_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_7_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_7_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_7_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_7_4"};

localparam string gather_rt_file_list_1_8[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_8_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_8_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_8_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_8_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_8_4"};

localparam string gather_rt_file_list_1_9[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_9_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_9_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_9_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_9_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_9_4"};

localparam string gather_rt_file_list_1_10[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_10_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_10_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_10_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_10_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_10_4"};

localparam string gather_rt_file_list_1_11[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_11_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_11_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_11_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_11_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_11_4"};

localparam string gather_rt_file_list_1_12[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_12_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_12_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_12_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_12_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_12_4"};

localparam string gather_rt_file_list_1_13[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_13_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_13_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_13_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_13_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_13_4"};

localparam string gather_rt_file_list_1_14[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_14_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_14_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_14_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_14_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_14_4"};

localparam string gather_rt_file_list_1_15[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_15_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_15_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_15_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_15_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_15_4"};

localparam string gather_rt_file_list_1_16[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_16_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_16_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_16_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_16_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_16_4"};

localparam string gather_rt_file_list_1_17[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_17_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_17_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_17_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_17_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_17_4"};

localparam string gather_rt_file_list_1_18[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_18_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_18_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_18_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_18_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_18_4"};

localparam string gather_rt_file_list_1_19[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_19_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_19_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_19_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_19_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_19_4"};

localparam string gather_rt_file_list_1_20[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_20_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_20_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_20_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_20_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_20_4"};

localparam string gather_rt_file_list_1_21[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_21_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_21_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_21_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_21_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_21_4"};

localparam string gather_rt_file_list_1_22[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_22_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_22_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_22_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_22_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_22_4"};

localparam string gather_rt_file_list_1_23[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_23_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_23_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_23_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_23_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_23_4"};

localparam string gather_rt_file_list_1_24[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_24_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_24_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_24_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_24_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_1_24_4"};

localparam string gather_rt_file_list_2_0[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_0_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_0_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_0_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_0_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_0_4"};

localparam string gather_rt_file_list_2_1[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_1_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_1_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_1_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_1_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_1_4"};

localparam string gather_rt_file_list_2_2[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_2_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_2_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_2_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_2_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_2_4"};

localparam string gather_rt_file_list_2_3[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_3_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_3_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_3_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_3_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_3_4"};

localparam string gather_rt_file_list_2_4[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_4_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_4_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_4_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_4_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_4_4"};

localparam string gather_rt_file_list_2_5[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_5_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_5_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_5_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_5_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_5_4"};

localparam string gather_rt_file_list_2_6[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_6_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_6_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_6_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_6_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_6_4"};

localparam string gather_rt_file_list_2_7[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_7_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_7_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_7_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_7_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_7_4"};

localparam string gather_rt_file_list_2_8[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_8_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_8_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_8_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_8_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_8_4"};

localparam string gather_rt_file_list_2_9[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_9_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_9_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_9_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_9_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_9_4"};

localparam string gather_rt_file_list_2_10[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_10_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_10_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_10_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_10_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_10_4"};

localparam string gather_rt_file_list_2_11[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_11_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_11_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_11_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_11_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_11_4"};

localparam string gather_rt_file_list_2_12[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_12_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_12_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_12_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_12_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_12_4"};

localparam string gather_rt_file_list_2_13[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_13_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_13_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_13_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_13_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_13_4"};

localparam string gather_rt_file_list_2_14[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_14_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_14_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_14_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_14_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_14_4"};

localparam string gather_rt_file_list_2_15[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_15_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_15_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_15_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_15_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_15_4"};

localparam string gather_rt_file_list_2_16[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_16_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_16_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_16_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_16_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_16_4"};

localparam string gather_rt_file_list_2_17[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_17_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_17_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_17_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_17_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_17_4"};

localparam string gather_rt_file_list_2_18[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_18_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_18_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_18_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_18_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_18_4"};

localparam string gather_rt_file_list_2_19[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_19_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_19_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_19_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_19_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_19_4"};

localparam string gather_rt_file_list_2_20[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_20_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_20_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_20_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_20_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_20_4"};

localparam string gather_rt_file_list_2_21[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_21_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_21_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_21_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_21_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_21_4"};

localparam string gather_rt_file_list_2_22[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_22_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_22_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_22_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_22_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_22_4"};

localparam string gather_rt_file_list_2_23[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_23_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_23_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_23_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_23_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_23_4"};

localparam string gather_rt_file_list_2_24[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_24_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_24_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_24_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_24_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_2_24_4"};

localparam string gather_rt_file_list_3_0[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_0_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_0_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_0_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_0_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_0_4"};

localparam string gather_rt_file_list_3_1[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_1_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_1_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_1_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_1_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_1_4"};

localparam string gather_rt_file_list_3_2[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_2_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_2_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_2_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_2_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_2_4"};

localparam string gather_rt_file_list_3_3[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_3_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_3_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_3_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_3_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_3_4"};

localparam string gather_rt_file_list_3_4[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_4_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_4_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_4_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_4_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_4_4"};

localparam string gather_rt_file_list_3_5[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_5_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_5_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_5_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_5_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_5_4"};

localparam string gather_rt_file_list_3_6[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_6_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_6_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_6_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_6_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_6_4"};

localparam string gather_rt_file_list_3_7[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_7_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_7_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_7_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_7_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_7_4"};

localparam string gather_rt_file_list_3_8[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_8_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_8_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_8_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_8_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_8_4"};

localparam string gather_rt_file_list_3_9[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_9_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_9_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_9_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_9_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_9_4"};

localparam string gather_rt_file_list_3_10[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_10_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_10_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_10_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_10_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_10_4"};

localparam string gather_rt_file_list_3_11[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_11_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_11_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_11_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_11_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_11_4"};

localparam string gather_rt_file_list_3_12[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_12_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_12_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_12_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_12_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_12_4"};

localparam string gather_rt_file_list_3_13[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_13_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_13_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_13_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_13_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_13_4"};

localparam string gather_rt_file_list_3_14[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_14_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_14_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_14_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_14_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_14_4"};

localparam string gather_rt_file_list_3_15[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_15_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_15_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_15_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_15_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_15_4"};

localparam string gather_rt_file_list_3_16[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_16_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_16_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_16_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_16_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_16_4"};

localparam string gather_rt_file_list_3_17[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_17_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_17_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_17_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_17_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_17_4"};

localparam string gather_rt_file_list_3_18[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_18_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_18_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_18_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_18_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_18_4"};

localparam string gather_rt_file_list_3_19[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_19_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_19_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_19_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_19_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_19_4"};

localparam string gather_rt_file_list_3_20[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_20_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_20_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_20_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_20_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_20_4"};

localparam string gather_rt_file_list_3_21[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_21_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_21_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_21_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_21_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_21_4"};

localparam string gather_rt_file_list_3_22[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_22_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_22_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_22_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_22_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_22_4"};

localparam string gather_rt_file_list_3_23[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_23_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_23_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_23_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_23_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_23_4"};

localparam string gather_rt_file_list_3_24[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_24_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_24_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_24_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_24_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_3_24_4"};

localparam string gather_rt_file_list_4_0[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_0_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_0_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_0_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_0_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_0_4"};

localparam string gather_rt_file_list_4_1[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_1_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_1_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_1_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_1_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_1_4"};

localparam string gather_rt_file_list_4_2[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_2_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_2_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_2_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_2_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_2_4"};

localparam string gather_rt_file_list_4_3[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_3_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_3_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_3_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_3_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_3_4"};

localparam string gather_rt_file_list_4_4[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_4_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_4_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_4_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_4_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_4_4"};

localparam string gather_rt_file_list_4_5[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_5_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_5_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_5_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_5_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_5_4"};

localparam string gather_rt_file_list_4_6[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_6_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_6_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_6_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_6_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_6_4"};

localparam string gather_rt_file_list_4_7[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_7_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_7_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_7_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_7_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_7_4"};

localparam string gather_rt_file_list_4_8[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_8_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_8_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_8_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_8_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_8_4"};

localparam string gather_rt_file_list_4_9[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_9_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_9_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_9_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_9_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_9_4"};

localparam string gather_rt_file_list_4_10[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_10_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_10_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_10_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_10_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_10_4"};

localparam string gather_rt_file_list_4_11[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_11_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_11_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_11_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_11_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_11_4"};

localparam string gather_rt_file_list_4_12[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_12_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_12_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_12_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_12_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_12_4"};

localparam string gather_rt_file_list_4_13[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_13_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_13_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_13_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_13_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_13_4"};

localparam string gather_rt_file_list_4_14[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_14_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_14_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_14_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_14_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_14_4"};

localparam string gather_rt_file_list_4_15[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_15_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_15_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_15_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_15_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_15_4"};

localparam string gather_rt_file_list_4_16[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_16_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_16_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_16_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_16_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_16_4"};

localparam string gather_rt_file_list_4_17[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_17_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_17_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_17_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_17_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_17_4"};

localparam string gather_rt_file_list_4_18[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_18_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_18_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_18_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_18_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_18_4"};

localparam string gather_rt_file_list_4_19[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_19_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_19_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_19_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_19_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_19_4"};

localparam string gather_rt_file_list_4_20[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_20_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_20_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_20_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_20_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_20_4"};

localparam string gather_rt_file_list_4_21[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_21_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_21_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_21_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_21_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_21_4"};

localparam string gather_rt_file_list_4_22[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_22_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_22_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_22_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_22_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_22_4"};

localparam string gather_rt_file_list_4_23[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_23_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_23_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_23_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_23_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_23_4"};

localparam string gather_rt_file_list_4_24[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_24_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_24_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_24_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_24_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_4_24_4"};

localparam string gather_rt_file_list_5_0[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_0_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_0_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_0_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_0_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_0_4"};

localparam string gather_rt_file_list_5_1[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_1_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_1_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_1_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_1_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_1_4"};

localparam string gather_rt_file_list_5_2[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_2_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_2_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_2_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_2_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_2_4"};

localparam string gather_rt_file_list_5_3[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_3_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_3_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_3_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_3_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_3_4"};

localparam string gather_rt_file_list_5_4[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_4_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_4_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_4_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_4_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_4_4"};

localparam string gather_rt_file_list_5_5[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_5_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_5_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_5_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_5_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_5_4"};

localparam string gather_rt_file_list_5_6[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_6_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_6_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_6_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_6_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_6_4"};

localparam string gather_rt_file_list_5_7[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_7_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_7_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_7_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_7_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_7_4"};

localparam string gather_rt_file_list_5_8[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_8_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_8_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_8_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_8_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_8_4"};

localparam string gather_rt_file_list_5_9[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_9_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_9_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_9_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_9_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_9_4"};

localparam string gather_rt_file_list_5_10[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_10_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_10_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_10_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_10_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_10_4"};

localparam string gather_rt_file_list_5_11[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_11_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_11_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_11_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_11_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_11_4"};

localparam string gather_rt_file_list_5_12[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_12_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_12_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_12_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_12_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_12_4"};

localparam string gather_rt_file_list_5_13[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_13_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_13_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_13_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_13_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_13_4"};

localparam string gather_rt_file_list_5_14[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_14_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_14_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_14_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_14_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_14_4"};

localparam string gather_rt_file_list_5_15[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_15_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_15_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_15_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_15_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_15_4"};

localparam string gather_rt_file_list_5_16[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_16_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_16_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_16_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_16_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_16_4"};

localparam string gather_rt_file_list_5_17[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_17_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_17_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_17_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_17_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_17_4"};

localparam string gather_rt_file_list_5_18[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_18_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_18_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_18_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_18_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_18_4"};

localparam string gather_rt_file_list_5_19[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_19_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_19_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_19_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_19_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_19_4"};

localparam string gather_rt_file_list_5_20[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_20_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_20_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_20_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_20_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_20_4"};

localparam string gather_rt_file_list_5_21[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_21_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_21_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_21_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_21_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_21_4"};

localparam string gather_rt_file_list_5_22[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_22_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_22_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_22_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_22_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_22_4"};

localparam string gather_rt_file_list_5_23[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_23_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_23_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_23_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_23_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_23_4"};

localparam string gather_rt_file_list_5_24[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_24_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_24_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_24_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_24_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_5_24_4"};

localparam string gather_rt_file_list_6_0[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_0_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_0_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_0_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_0_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_0_4"};

localparam string gather_rt_file_list_6_1[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_1_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_1_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_1_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_1_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_1_4"};

localparam string gather_rt_file_list_6_2[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_2_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_2_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_2_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_2_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_2_4"};

localparam string gather_rt_file_list_6_3[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_3_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_3_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_3_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_3_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_3_4"};

localparam string gather_rt_file_list_6_4[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_4_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_4_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_4_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_4_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_4_4"};

localparam string gather_rt_file_list_6_5[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_5_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_5_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_5_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_5_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_5_4"};

localparam string gather_rt_file_list_6_6[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_6_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_6_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_6_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_6_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_6_4"};

localparam string gather_rt_file_list_6_7[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_7_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_7_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_7_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_7_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_7_4"};

localparam string gather_rt_file_list_6_8[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_8_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_8_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_8_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_8_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_8_4"};

localparam string gather_rt_file_list_6_9[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_9_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_9_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_9_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_9_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_9_4"};

localparam string gather_rt_file_list_6_10[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_10_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_10_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_10_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_10_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_10_4"};

localparam string gather_rt_file_list_6_11[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_11_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_11_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_11_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_11_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_11_4"};

localparam string gather_rt_file_list_6_12[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_12_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_12_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_12_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_12_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_12_4"};

localparam string gather_rt_file_list_6_13[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_13_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_13_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_13_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_13_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_13_4"};

localparam string gather_rt_file_list_6_14[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_14_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_14_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_14_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_14_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_14_4"};

localparam string gather_rt_file_list_6_15[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_15_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_15_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_15_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_15_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_15_4"};

localparam string gather_rt_file_list_6_16[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_16_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_16_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_16_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_16_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_16_4"};

localparam string gather_rt_file_list_6_17[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_17_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_17_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_17_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_17_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_17_4"};

localparam string gather_rt_file_list_6_18[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_18_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_18_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_18_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_18_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_18_4"};

localparam string gather_rt_file_list_6_19[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_19_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_19_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_19_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_19_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_19_4"};

localparam string gather_rt_file_list_6_20[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_20_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_20_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_20_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_20_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_20_4"};

localparam string gather_rt_file_list_6_21[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_21_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_21_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_21_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_21_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_21_4"};

localparam string gather_rt_file_list_6_22[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_22_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_22_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_22_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_22_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_22_4"};

localparam string gather_rt_file_list_6_23[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_23_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_23_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_23_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_23_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_23_4"};

localparam string gather_rt_file_list_6_24[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_24_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_24_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_24_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_24_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_6_24_4"};

localparam string gather_rt_file_list_7_0[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_0_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_0_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_0_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_0_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_0_4"};

localparam string gather_rt_file_list_7_1[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_1_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_1_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_1_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_1_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_1_4"};

localparam string gather_rt_file_list_7_2[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_2_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_2_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_2_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_2_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_2_4"};

localparam string gather_rt_file_list_7_3[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_3_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_3_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_3_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_3_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_3_4"};

localparam string gather_rt_file_list_7_4[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_4_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_4_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_4_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_4_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_4_4"};

localparam string gather_rt_file_list_7_5[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_5_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_5_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_5_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_5_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_5_4"};

localparam string gather_rt_file_list_7_6[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_6_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_6_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_6_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_6_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_6_4"};

localparam string gather_rt_file_list_7_7[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_7_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_7_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_7_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_7_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_7_4"};

localparam string gather_rt_file_list_7_8[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_8_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_8_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_8_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_8_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_8_4"};

localparam string gather_rt_file_list_7_9[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_9_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_9_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_9_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_9_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_9_4"};

localparam string gather_rt_file_list_7_10[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_10_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_10_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_10_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_10_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_10_4"};

localparam string gather_rt_file_list_7_11[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_11_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_11_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_11_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_11_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_11_4"};

localparam string gather_rt_file_list_7_12[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_12_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_12_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_12_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_12_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_12_4"};

localparam string gather_rt_file_list_7_13[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_13_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_13_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_13_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_13_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_13_4"};

localparam string gather_rt_file_list_7_14[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_14_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_14_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_14_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_14_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_14_4"};

localparam string gather_rt_file_list_7_15[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_15_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_15_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_15_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_15_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_15_4"};

localparam string gather_rt_file_list_7_16[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_16_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_16_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_16_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_16_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_16_4"};

localparam string gather_rt_file_list_7_17[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_17_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_17_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_17_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_17_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_17_4"};

localparam string gather_rt_file_list_7_18[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_18_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_18_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_18_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_18_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_18_4"};

localparam string gather_rt_file_list_7_19[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_19_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_19_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_19_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_19_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_19_4"};

localparam string gather_rt_file_list_7_20[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_20_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_20_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_20_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_20_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_20_4"};

localparam string gather_rt_file_list_7_21[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_21_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_21_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_21_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_21_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_21_4"};

localparam string gather_rt_file_list_7_22[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_22_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_22_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_22_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_22_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_22_4"};

localparam string gather_rt_file_list_7_23[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_23_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_23_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_23_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_23_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_23_4"};

localparam string gather_rt_file_list_7_24[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_24_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_24_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_24_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_24_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_7_24_4"};

localparam string gather_rt_file_list_8_0[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_0_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_0_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_0_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_0_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_0_4"};

localparam string gather_rt_file_list_8_1[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_1_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_1_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_1_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_1_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_1_4"};

localparam string gather_rt_file_list_8_2[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_2_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_2_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_2_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_2_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_2_4"};

localparam string gather_rt_file_list_8_3[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_3_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_3_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_3_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_3_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_3_4"};

localparam string gather_rt_file_list_8_4[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_4_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_4_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_4_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_4_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_4_4"};

localparam string gather_rt_file_list_8_5[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_5_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_5_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_5_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_5_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_5_4"};

localparam string gather_rt_file_list_8_6[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_6_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_6_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_6_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_6_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_6_4"};

localparam string gather_rt_file_list_8_7[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_7_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_7_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_7_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_7_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_7_4"};

localparam string gather_rt_file_list_8_8[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_8_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_8_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_8_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_8_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_8_4"};

localparam string gather_rt_file_list_8_9[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_9_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_9_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_9_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_9_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_9_4"};

localparam string gather_rt_file_list_8_10[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_10_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_10_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_10_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_10_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_10_4"};

localparam string gather_rt_file_list_8_11[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_11_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_11_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_11_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_11_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_11_4"};

localparam string gather_rt_file_list_8_12[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_12_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_12_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_12_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_12_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_12_4"};

localparam string gather_rt_file_list_8_13[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_13_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_13_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_13_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_13_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_13_4"};

localparam string gather_rt_file_list_8_14[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_14_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_14_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_14_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_14_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_14_4"};

localparam string gather_rt_file_list_8_15[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_15_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_15_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_15_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_15_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_15_4"};

localparam string gather_rt_file_list_8_16[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_16_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_16_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_16_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_16_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_16_4"};

localparam string gather_rt_file_list_8_17[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_17_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_17_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_17_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_17_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_17_4"};

localparam string gather_rt_file_list_8_18[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_18_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_18_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_18_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_18_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_18_4"};

localparam string gather_rt_file_list_8_19[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_19_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_19_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_19_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_19_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_19_4"};

localparam string gather_rt_file_list_8_20[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_20_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_20_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_20_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_20_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_20_4"};

localparam string gather_rt_file_list_8_21[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_21_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_21_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_21_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_21_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_21_4"};

localparam string gather_rt_file_list_8_22[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_22_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_22_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_22_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_22_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_22_4"};

localparam string gather_rt_file_list_8_23[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_23_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_23_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_23_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_23_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_23_4"};

localparam string gather_rt_file_list_8_24[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_24_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_24_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_24_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_24_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_8_24_4"};

localparam string gather_rt_file_list_9_0[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_0_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_0_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_0_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_0_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_0_4"};

localparam string gather_rt_file_list_9_1[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_1_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_1_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_1_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_1_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_1_4"};

localparam string gather_rt_file_list_9_2[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_2_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_2_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_2_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_2_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_2_4"};

localparam string gather_rt_file_list_9_3[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_3_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_3_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_3_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_3_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_3_4"};

localparam string gather_rt_file_list_9_4[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_4_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_4_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_4_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_4_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_4_4"};

localparam string gather_rt_file_list_9_5[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_5_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_5_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_5_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_5_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_5_4"};

localparam string gather_rt_file_list_9_6[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_6_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_6_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_6_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_6_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_6_4"};

localparam string gather_rt_file_list_9_7[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_7_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_7_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_7_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_7_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_7_4"};

localparam string gather_rt_file_list_9_8[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_8_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_8_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_8_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_8_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_8_4"};

localparam string gather_rt_file_list_9_9[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_9_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_9_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_9_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_9_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_9_4"};

localparam string gather_rt_file_list_9_10[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_10_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_10_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_10_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_10_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_10_4"};

localparam string gather_rt_file_list_9_11[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_11_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_11_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_11_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_11_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_11_4"};

localparam string gather_rt_file_list_9_12[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_12_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_12_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_12_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_12_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_12_4"};

localparam string gather_rt_file_list_9_13[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_13_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_13_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_13_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_13_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_13_4"};

localparam string gather_rt_file_list_9_14[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_14_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_14_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_14_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_14_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_14_4"};

localparam string gather_rt_file_list_9_15[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_15_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_15_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_15_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_15_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_15_4"};

localparam string gather_rt_file_list_9_16[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_16_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_16_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_16_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_16_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_16_4"};

localparam string gather_rt_file_list_9_17[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_17_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_17_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_17_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_17_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_17_4"};

localparam string gather_rt_file_list_9_18[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_18_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_18_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_18_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_18_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_18_4"};

localparam string gather_rt_file_list_9_19[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_19_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_19_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_19_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_19_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_19_4"};

localparam string gather_rt_file_list_9_20[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_20_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_20_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_20_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_20_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_20_4"};

localparam string gather_rt_file_list_9_21[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_21_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_21_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_21_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_21_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_21_4"};

localparam string gather_rt_file_list_9_22[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_22_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_22_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_22_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_22_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_22_4"};

localparam string gather_rt_file_list_9_23[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_23_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_23_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_23_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_23_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_23_4"};

localparam string gather_rt_file_list_9_24[`CN] = '{"/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_24_0","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_24_1","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_24_2","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_24_3","/mnt/c/git/nvcim-comm/network/config/routing_tables/gather_9_24_4"};

`endif
