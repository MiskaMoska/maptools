`include "params.svh"
`include "network_config.svh"

module system (
    input       wire                            clk,
    input       wire                            rstn,

    input       wire        [`DW-1:0]           data_i_stab,
    input       wire                            valid_i_stab,
    output      wire                            ready_o_stab,

    output      wire        [`DW-1:0]           data_o_flee0,
    output      wire                            valid_o_flee0,
    input       wire                            ready_i_flee0,

    output      wire        [`DW-1:0]           data_o_flee1,
    output      wire                            valid_o_flee1,
    input       wire                            ready_i_flee1  
);

wire [`DW-1:0] cast_data_pe_2_nw[`NOC_WIDTH][`NOC_HEIGHT], merge_data_pe_2_nw[`NOC_WIDTH][`NOC_HEIGHT], cast_data_nw_2_pe[`NOC_WIDTH][`NOC_HEIGHT], merge_data_nw_2_pe[`NOC_WIDTH][`NOC_HEIGHT];
wire  cast_valid_pe_2_nw[`NOC_WIDTH][`NOC_HEIGHT], merge_valid_pe_2_nw[`NOC_WIDTH][`NOC_HEIGHT], cast_valid_nw_2_pe[`NOC_WIDTH][`NOC_HEIGHT], merge_valid_nw_2_pe[`NOC_WIDTH][`NOC_HEIGHT];
wire  cast_ready_pe_2_nw[`NOC_WIDTH][`NOC_HEIGHT], merge_ready_pe_2_nw[`NOC_WIDTH][`NOC_HEIGHT], cast_ready_nw_2_pe[`NOC_WIDTH][`NOC_HEIGHT], merge_ready_nw_2_pe[`NOC_WIDTH][`NOC_HEIGHT];

network nw(
    .clk                                                  (clk),
    .rstn                                                 (rstn),
    .data_i_stab                                          (data_i_stab),
    .valid_i_stab                                         (valid_i_stab),
    .ready_o_stab                                         (ready_o_stab),
    .data_o_flee0                                         (data_o_flee0),
    .valid_o_flee0                                        (valid_o_flee0),
    .ready_i_flee0                                        (ready_i_flee0),
    .data_o_flee1                                         (data_o_flee1),
    .valid_o_flee1                                        (valid_o_flee1),
    .ready_i_flee1                                        (ready_i_flee1),
    .cast_data_i                                          (cast_data_pe_2_nw),
    .cast_valid_i                                         (cast_valid_pe_2_nw),
    .cast_ready_o                                         (cast_ready_nw_2_pe),
    .cast_data_o                                          (cast_data_nw_2_pe),
    .cast_valid_o                                         (cast_valid_nw_2_pe),
    .cast_ready_i                                         (cast_ready_pe_2_nw),
    .merge_data_i                                         (merge_data_pe_2_nw),
    .merge_valid_i                                        (merge_valid_pe_2_nw),
    .merge_ready_o                                        (merge_ready_nw_2_pe),
    .merge_data_o                                         (merge_data_nw_2_pe),
    .merge_valid_o                                        (merge_valid_nw_2_pe),
    .merge_ready_i                                        (merge_ready_pe_2_nw)
);

virtual_pe #(
    .isCaster                    (isCaster_0_0)
)vpe_0_0(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[0][0]),
    .cast_valid_i                (cast_valid_nw_2_pe[0][0]),
    .cast_ready_o                (cast_ready_pe_2_nw[0][0]),
    .cast_data_o                 (cast_data_pe_2_nw[0][0]),
    .cast_valid_o                (cast_valid_pe_2_nw[0][0]),
    .cast_ready_i                (cast_ready_nw_2_pe[0][0]),
    .merge_data_i                (merge_data_nw_2_pe[0][0]),
    .merge_valid_i               (merge_valid_nw_2_pe[0][0]),
    .merge_ready_o               (merge_ready_pe_2_nw[0][0]),
    .merge_data_o                (merge_data_pe_2_nw[0][0]),
    .merge_valid_o               (merge_valid_pe_2_nw[0][0]),
    .merge_ready_i               (merge_ready_nw_2_pe[0][0])
);


virtual_pe #(
    .isCaster                    (isCaster_0_1)
)vpe_0_1(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[0][1]),
    .cast_valid_i                (cast_valid_nw_2_pe[0][1]),
    .cast_ready_o                (cast_ready_pe_2_nw[0][1]),
    .cast_data_o                 (cast_data_pe_2_nw[0][1]),
    .cast_valid_o                (cast_valid_pe_2_nw[0][1]),
    .cast_ready_i                (cast_ready_nw_2_pe[0][1]),
    .merge_data_i                (merge_data_nw_2_pe[0][1]),
    .merge_valid_i               (merge_valid_nw_2_pe[0][1]),
    .merge_ready_o               (merge_ready_pe_2_nw[0][1]),
    .merge_data_o                (merge_data_pe_2_nw[0][1]),
    .merge_valid_o               (merge_valid_pe_2_nw[0][1]),
    .merge_ready_i               (merge_ready_nw_2_pe[0][1])
);


virtual_pe #(
    .isCaster                    (isCaster_0_2)
)vpe_0_2(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[0][2]),
    .cast_valid_i                (cast_valid_nw_2_pe[0][2]),
    .cast_ready_o                (cast_ready_pe_2_nw[0][2]),
    .cast_data_o                 (cast_data_pe_2_nw[0][2]),
    .cast_valid_o                (cast_valid_pe_2_nw[0][2]),
    .cast_ready_i                (cast_ready_nw_2_pe[0][2]),
    .merge_data_i                (merge_data_nw_2_pe[0][2]),
    .merge_valid_i               (merge_valid_nw_2_pe[0][2]),
    .merge_ready_o               (merge_ready_pe_2_nw[0][2]),
    .merge_data_o                (merge_data_pe_2_nw[0][2]),
    .merge_valid_o               (merge_valid_pe_2_nw[0][2]),
    .merge_ready_i               (merge_ready_nw_2_pe[0][2])
);


virtual_pe #(
    .isCaster                    (isCaster_0_3)
)vpe_0_3(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[0][3]),
    .cast_valid_i                (cast_valid_nw_2_pe[0][3]),
    .cast_ready_o                (cast_ready_pe_2_nw[0][3]),
    .cast_data_o                 (cast_data_pe_2_nw[0][3]),
    .cast_valid_o                (cast_valid_pe_2_nw[0][3]),
    .cast_ready_i                (cast_ready_nw_2_pe[0][3]),
    .merge_data_i                (merge_data_nw_2_pe[0][3]),
    .merge_valid_i               (merge_valid_nw_2_pe[0][3]),
    .merge_ready_o               (merge_ready_pe_2_nw[0][3]),
    .merge_data_o                (merge_data_pe_2_nw[0][3]),
    .merge_valid_o               (merge_valid_pe_2_nw[0][3]),
    .merge_ready_i               (merge_ready_nw_2_pe[0][3])
);


virtual_pe #(
    .isCaster                    (isCaster_0_4)
)vpe_0_4(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[0][4]),
    .cast_valid_i                (cast_valid_nw_2_pe[0][4]),
    .cast_ready_o                (cast_ready_pe_2_nw[0][4]),
    .cast_data_o                 (cast_data_pe_2_nw[0][4]),
    .cast_valid_o                (cast_valid_pe_2_nw[0][4]),
    .cast_ready_i                (cast_ready_nw_2_pe[0][4]),
    .merge_data_i                (merge_data_nw_2_pe[0][4]),
    .merge_valid_i               (merge_valid_nw_2_pe[0][4]),
    .merge_ready_o               (merge_ready_pe_2_nw[0][4]),
    .merge_data_o                (merge_data_pe_2_nw[0][4]),
    .merge_valid_o               (merge_valid_pe_2_nw[0][4]),
    .merge_ready_i               (merge_ready_nw_2_pe[0][4])
);


virtual_pe #(
    .isCaster                    (isCaster_0_5)
)vpe_0_5(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[0][5]),
    .cast_valid_i                (cast_valid_nw_2_pe[0][5]),
    .cast_ready_o                (cast_ready_pe_2_nw[0][5]),
    .cast_data_o                 (cast_data_pe_2_nw[0][5]),
    .cast_valid_o                (cast_valid_pe_2_nw[0][5]),
    .cast_ready_i                (cast_ready_nw_2_pe[0][5]),
    .merge_data_i                (merge_data_nw_2_pe[0][5]),
    .merge_valid_i               (merge_valid_nw_2_pe[0][5]),
    .merge_ready_o               (merge_ready_pe_2_nw[0][5]),
    .merge_data_o                (merge_data_pe_2_nw[0][5]),
    .merge_valid_o               (merge_valid_pe_2_nw[0][5]),
    .merge_ready_i               (merge_ready_nw_2_pe[0][5])
);


virtual_pe #(
    .isCaster                    (isCaster_0_6)
)vpe_0_6(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[0][6]),
    .cast_valid_i                (cast_valid_nw_2_pe[0][6]),
    .cast_ready_o                (cast_ready_pe_2_nw[0][6]),
    .cast_data_o                 (cast_data_pe_2_nw[0][6]),
    .cast_valid_o                (cast_valid_pe_2_nw[0][6]),
    .cast_ready_i                (cast_ready_nw_2_pe[0][6]),
    .merge_data_i                (merge_data_nw_2_pe[0][6]),
    .merge_valid_i               (merge_valid_nw_2_pe[0][6]),
    .merge_ready_o               (merge_ready_pe_2_nw[0][6]),
    .merge_data_o                (merge_data_pe_2_nw[0][6]),
    .merge_valid_o               (merge_valid_pe_2_nw[0][6]),
    .merge_ready_i               (merge_ready_nw_2_pe[0][6])
);


virtual_pe #(
    .isCaster                    (isCaster_0_7)
)vpe_0_7(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[0][7]),
    .cast_valid_i                (cast_valid_nw_2_pe[0][7]),
    .cast_ready_o                (cast_ready_pe_2_nw[0][7]),
    .cast_data_o                 (cast_data_pe_2_nw[0][7]),
    .cast_valid_o                (cast_valid_pe_2_nw[0][7]),
    .cast_ready_i                (cast_ready_nw_2_pe[0][7]),
    .merge_data_i                (merge_data_nw_2_pe[0][7]),
    .merge_valid_i               (merge_valid_nw_2_pe[0][7]),
    .merge_ready_o               (merge_ready_pe_2_nw[0][7]),
    .merge_data_o                (merge_data_pe_2_nw[0][7]),
    .merge_valid_o               (merge_valid_pe_2_nw[0][7]),
    .merge_ready_i               (merge_ready_nw_2_pe[0][7])
);


virtual_pe #(
    .isCaster                    (isCaster_1_0)
)vpe_1_0(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[1][0]),
    .cast_valid_i                (cast_valid_nw_2_pe[1][0]),
    .cast_ready_o                (cast_ready_pe_2_nw[1][0]),
    .cast_data_o                 (cast_data_pe_2_nw[1][0]),
    .cast_valid_o                (cast_valid_pe_2_nw[1][0]),
    .cast_ready_i                (cast_ready_nw_2_pe[1][0]),
    .merge_data_i                (merge_data_nw_2_pe[1][0]),
    .merge_valid_i               (merge_valid_nw_2_pe[1][0]),
    .merge_ready_o               (merge_ready_pe_2_nw[1][0]),
    .merge_data_o                (merge_data_pe_2_nw[1][0]),
    .merge_valid_o               (merge_valid_pe_2_nw[1][0]),
    .merge_ready_i               (merge_ready_nw_2_pe[1][0])
);


virtual_pe #(
    .isCaster                    (isCaster_1_1)
)vpe_1_1(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[1][1]),
    .cast_valid_i                (cast_valid_nw_2_pe[1][1]),
    .cast_ready_o                (cast_ready_pe_2_nw[1][1]),
    .cast_data_o                 (cast_data_pe_2_nw[1][1]),
    .cast_valid_o                (cast_valid_pe_2_nw[1][1]),
    .cast_ready_i                (cast_ready_nw_2_pe[1][1]),
    .merge_data_i                (merge_data_nw_2_pe[1][1]),
    .merge_valid_i               (merge_valid_nw_2_pe[1][1]),
    .merge_ready_o               (merge_ready_pe_2_nw[1][1]),
    .merge_data_o                (merge_data_pe_2_nw[1][1]),
    .merge_valid_o               (merge_valid_pe_2_nw[1][1]),
    .merge_ready_i               (merge_ready_nw_2_pe[1][1])
);


virtual_pe #(
    .isCaster                    (isCaster_1_2)
)vpe_1_2(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[1][2]),
    .cast_valid_i                (cast_valid_nw_2_pe[1][2]),
    .cast_ready_o                (cast_ready_pe_2_nw[1][2]),
    .cast_data_o                 (cast_data_pe_2_nw[1][2]),
    .cast_valid_o                (cast_valid_pe_2_nw[1][2]),
    .cast_ready_i                (cast_ready_nw_2_pe[1][2]),
    .merge_data_i                (merge_data_nw_2_pe[1][2]),
    .merge_valid_i               (merge_valid_nw_2_pe[1][2]),
    .merge_ready_o               (merge_ready_pe_2_nw[1][2]),
    .merge_data_o                (merge_data_pe_2_nw[1][2]),
    .merge_valid_o               (merge_valid_pe_2_nw[1][2]),
    .merge_ready_i               (merge_ready_nw_2_pe[1][2])
);


virtual_pe #(
    .isCaster                    (isCaster_1_3)
)vpe_1_3(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[1][3]),
    .cast_valid_i                (cast_valid_nw_2_pe[1][3]),
    .cast_ready_o                (cast_ready_pe_2_nw[1][3]),
    .cast_data_o                 (cast_data_pe_2_nw[1][3]),
    .cast_valid_o                (cast_valid_pe_2_nw[1][3]),
    .cast_ready_i                (cast_ready_nw_2_pe[1][3]),
    .merge_data_i                (merge_data_nw_2_pe[1][3]),
    .merge_valid_i               (merge_valid_nw_2_pe[1][3]),
    .merge_ready_o               (merge_ready_pe_2_nw[1][3]),
    .merge_data_o                (merge_data_pe_2_nw[1][3]),
    .merge_valid_o               (merge_valid_pe_2_nw[1][3]),
    .merge_ready_i               (merge_ready_nw_2_pe[1][3])
);


virtual_pe #(
    .isCaster                    (isCaster_1_4)
)vpe_1_4(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[1][4]),
    .cast_valid_i                (cast_valid_nw_2_pe[1][4]),
    .cast_ready_o                (cast_ready_pe_2_nw[1][4]),
    .cast_data_o                 (cast_data_pe_2_nw[1][4]),
    .cast_valid_o                (cast_valid_pe_2_nw[1][4]),
    .cast_ready_i                (cast_ready_nw_2_pe[1][4]),
    .merge_data_i                (merge_data_nw_2_pe[1][4]),
    .merge_valid_i               (merge_valid_nw_2_pe[1][4]),
    .merge_ready_o               (merge_ready_pe_2_nw[1][4]),
    .merge_data_o                (merge_data_pe_2_nw[1][4]),
    .merge_valid_o               (merge_valid_pe_2_nw[1][4]),
    .merge_ready_i               (merge_ready_nw_2_pe[1][4])
);


virtual_pe #(
    .isCaster                    (isCaster_1_5)
)vpe_1_5(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[1][5]),
    .cast_valid_i                (cast_valid_nw_2_pe[1][5]),
    .cast_ready_o                (cast_ready_pe_2_nw[1][5]),
    .cast_data_o                 (cast_data_pe_2_nw[1][5]),
    .cast_valid_o                (cast_valid_pe_2_nw[1][5]),
    .cast_ready_i                (cast_ready_nw_2_pe[1][5]),
    .merge_data_i                (merge_data_nw_2_pe[1][5]),
    .merge_valid_i               (merge_valid_nw_2_pe[1][5]),
    .merge_ready_o               (merge_ready_pe_2_nw[1][5]),
    .merge_data_o                (merge_data_pe_2_nw[1][5]),
    .merge_valid_o               (merge_valid_pe_2_nw[1][5]),
    .merge_ready_i               (merge_ready_nw_2_pe[1][5])
);


virtual_pe #(
    .isCaster                    (isCaster_1_6)
)vpe_1_6(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[1][6]),
    .cast_valid_i                (cast_valid_nw_2_pe[1][6]),
    .cast_ready_o                (cast_ready_pe_2_nw[1][6]),
    .cast_data_o                 (cast_data_pe_2_nw[1][6]),
    .cast_valid_o                (cast_valid_pe_2_nw[1][6]),
    .cast_ready_i                (cast_ready_nw_2_pe[1][6]),
    .merge_data_i                (merge_data_nw_2_pe[1][6]),
    .merge_valid_i               (merge_valid_nw_2_pe[1][6]),
    .merge_ready_o               (merge_ready_pe_2_nw[1][6]),
    .merge_data_o                (merge_data_pe_2_nw[1][6]),
    .merge_valid_o               (merge_valid_pe_2_nw[1][6]),
    .merge_ready_i               (merge_ready_nw_2_pe[1][6])
);


virtual_pe #(
    .isCaster                    (isCaster_1_7)
)vpe_1_7(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[1][7]),
    .cast_valid_i                (cast_valid_nw_2_pe[1][7]),
    .cast_ready_o                (cast_ready_pe_2_nw[1][7]),
    .cast_data_o                 (cast_data_pe_2_nw[1][7]),
    .cast_valid_o                (cast_valid_pe_2_nw[1][7]),
    .cast_ready_i                (cast_ready_nw_2_pe[1][7]),
    .merge_data_i                (merge_data_nw_2_pe[1][7]),
    .merge_valid_i               (merge_valid_nw_2_pe[1][7]),
    .merge_ready_o               (merge_ready_pe_2_nw[1][7]),
    .merge_data_o                (merge_data_pe_2_nw[1][7]),
    .merge_valid_o               (merge_valid_pe_2_nw[1][7]),
    .merge_ready_i               (merge_ready_nw_2_pe[1][7])
);


virtual_pe #(
    .isCaster                    (isCaster_2_0)
)vpe_2_0(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[2][0]),
    .cast_valid_i                (cast_valid_nw_2_pe[2][0]),
    .cast_ready_o                (cast_ready_pe_2_nw[2][0]),
    .cast_data_o                 (cast_data_pe_2_nw[2][0]),
    .cast_valid_o                (cast_valid_pe_2_nw[2][0]),
    .cast_ready_i                (cast_ready_nw_2_pe[2][0]),
    .merge_data_i                (merge_data_nw_2_pe[2][0]),
    .merge_valid_i               (merge_valid_nw_2_pe[2][0]),
    .merge_ready_o               (merge_ready_pe_2_nw[2][0]),
    .merge_data_o                (merge_data_pe_2_nw[2][0]),
    .merge_valid_o               (merge_valid_pe_2_nw[2][0]),
    .merge_ready_i               (merge_ready_nw_2_pe[2][0])
);


virtual_pe #(
    .isCaster                    (isCaster_2_1)
)vpe_2_1(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[2][1]),
    .cast_valid_i                (cast_valid_nw_2_pe[2][1]),
    .cast_ready_o                (cast_ready_pe_2_nw[2][1]),
    .cast_data_o                 (cast_data_pe_2_nw[2][1]),
    .cast_valid_o                (cast_valid_pe_2_nw[2][1]),
    .cast_ready_i                (cast_ready_nw_2_pe[2][1]),
    .merge_data_i                (merge_data_nw_2_pe[2][1]),
    .merge_valid_i               (merge_valid_nw_2_pe[2][1]),
    .merge_ready_o               (merge_ready_pe_2_nw[2][1]),
    .merge_data_o                (merge_data_pe_2_nw[2][1]),
    .merge_valid_o               (merge_valid_pe_2_nw[2][1]),
    .merge_ready_i               (merge_ready_nw_2_pe[2][1])
);


virtual_pe #(
    .isCaster                    (isCaster_2_2)
)vpe_2_2(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[2][2]),
    .cast_valid_i                (cast_valid_nw_2_pe[2][2]),
    .cast_ready_o                (cast_ready_pe_2_nw[2][2]),
    .cast_data_o                 (cast_data_pe_2_nw[2][2]),
    .cast_valid_o                (cast_valid_pe_2_nw[2][2]),
    .cast_ready_i                (cast_ready_nw_2_pe[2][2]),
    .merge_data_i                (merge_data_nw_2_pe[2][2]),
    .merge_valid_i               (merge_valid_nw_2_pe[2][2]),
    .merge_ready_o               (merge_ready_pe_2_nw[2][2]),
    .merge_data_o                (merge_data_pe_2_nw[2][2]),
    .merge_valid_o               (merge_valid_pe_2_nw[2][2]),
    .merge_ready_i               (merge_ready_nw_2_pe[2][2])
);


virtual_pe #(
    .isCaster                    (isCaster_2_3)
)vpe_2_3(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[2][3]),
    .cast_valid_i                (cast_valid_nw_2_pe[2][3]),
    .cast_ready_o                (cast_ready_pe_2_nw[2][3]),
    .cast_data_o                 (cast_data_pe_2_nw[2][3]),
    .cast_valid_o                (cast_valid_pe_2_nw[2][3]),
    .cast_ready_i                (cast_ready_nw_2_pe[2][3]),
    .merge_data_i                (merge_data_nw_2_pe[2][3]),
    .merge_valid_i               (merge_valid_nw_2_pe[2][3]),
    .merge_ready_o               (merge_ready_pe_2_nw[2][3]),
    .merge_data_o                (merge_data_pe_2_nw[2][3]),
    .merge_valid_o               (merge_valid_pe_2_nw[2][3]),
    .merge_ready_i               (merge_ready_nw_2_pe[2][3])
);


virtual_pe #(
    .isCaster                    (isCaster_2_4)
)vpe_2_4(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[2][4]),
    .cast_valid_i                (cast_valid_nw_2_pe[2][4]),
    .cast_ready_o                (cast_ready_pe_2_nw[2][4]),
    .cast_data_o                 (cast_data_pe_2_nw[2][4]),
    .cast_valid_o                (cast_valid_pe_2_nw[2][4]),
    .cast_ready_i                (cast_ready_nw_2_pe[2][4]),
    .merge_data_i                (merge_data_nw_2_pe[2][4]),
    .merge_valid_i               (merge_valid_nw_2_pe[2][4]),
    .merge_ready_o               (merge_ready_pe_2_nw[2][4]),
    .merge_data_o                (merge_data_pe_2_nw[2][4]),
    .merge_valid_o               (merge_valid_pe_2_nw[2][4]),
    .merge_ready_i               (merge_ready_nw_2_pe[2][4])
);


virtual_pe #(
    .isCaster                    (isCaster_2_5)
)vpe_2_5(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[2][5]),
    .cast_valid_i                (cast_valid_nw_2_pe[2][5]),
    .cast_ready_o                (cast_ready_pe_2_nw[2][5]),
    .cast_data_o                 (cast_data_pe_2_nw[2][5]),
    .cast_valid_o                (cast_valid_pe_2_nw[2][5]),
    .cast_ready_i                (cast_ready_nw_2_pe[2][5]),
    .merge_data_i                (merge_data_nw_2_pe[2][5]),
    .merge_valid_i               (merge_valid_nw_2_pe[2][5]),
    .merge_ready_o               (merge_ready_pe_2_nw[2][5]),
    .merge_data_o                (merge_data_pe_2_nw[2][5]),
    .merge_valid_o               (merge_valid_pe_2_nw[2][5]),
    .merge_ready_i               (merge_ready_nw_2_pe[2][5])
);


virtual_pe #(
    .isCaster                    (isCaster_2_6)
)vpe_2_6(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[2][6]),
    .cast_valid_i                (cast_valid_nw_2_pe[2][6]),
    .cast_ready_o                (cast_ready_pe_2_nw[2][6]),
    .cast_data_o                 (cast_data_pe_2_nw[2][6]),
    .cast_valid_o                (cast_valid_pe_2_nw[2][6]),
    .cast_ready_i                (cast_ready_nw_2_pe[2][6]),
    .merge_data_i                (merge_data_nw_2_pe[2][6]),
    .merge_valid_i               (merge_valid_nw_2_pe[2][6]),
    .merge_ready_o               (merge_ready_pe_2_nw[2][6]),
    .merge_data_o                (merge_data_pe_2_nw[2][6]),
    .merge_valid_o               (merge_valid_pe_2_nw[2][6]),
    .merge_ready_i               (merge_ready_nw_2_pe[2][6])
);


virtual_pe #(
    .isCaster                    (isCaster_2_7)
)vpe_2_7(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[2][7]),
    .cast_valid_i                (cast_valid_nw_2_pe[2][7]),
    .cast_ready_o                (cast_ready_pe_2_nw[2][7]),
    .cast_data_o                 (cast_data_pe_2_nw[2][7]),
    .cast_valid_o                (cast_valid_pe_2_nw[2][7]),
    .cast_ready_i                (cast_ready_nw_2_pe[2][7]),
    .merge_data_i                (merge_data_nw_2_pe[2][7]),
    .merge_valid_i               (merge_valid_nw_2_pe[2][7]),
    .merge_ready_o               (merge_ready_pe_2_nw[2][7]),
    .merge_data_o                (merge_data_pe_2_nw[2][7]),
    .merge_valid_o               (merge_valid_pe_2_nw[2][7]),
    .merge_ready_i               (merge_ready_nw_2_pe[2][7])
);


virtual_pe #(
    .isCaster                    (isCaster_3_0)
)vpe_3_0(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[3][0]),
    .cast_valid_i                (cast_valid_nw_2_pe[3][0]),
    .cast_ready_o                (cast_ready_pe_2_nw[3][0]),
    .cast_data_o                 (cast_data_pe_2_nw[3][0]),
    .cast_valid_o                (cast_valid_pe_2_nw[3][0]),
    .cast_ready_i                (cast_ready_nw_2_pe[3][0]),
    .merge_data_i                (merge_data_nw_2_pe[3][0]),
    .merge_valid_i               (merge_valid_nw_2_pe[3][0]),
    .merge_ready_o               (merge_ready_pe_2_nw[3][0]),
    .merge_data_o                (merge_data_pe_2_nw[3][0]),
    .merge_valid_o               (merge_valid_pe_2_nw[3][0]),
    .merge_ready_i               (merge_ready_nw_2_pe[3][0])
);


virtual_pe #(
    .isCaster                    (isCaster_3_1)
)vpe_3_1(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[3][1]),
    .cast_valid_i                (cast_valid_nw_2_pe[3][1]),
    .cast_ready_o                (cast_ready_pe_2_nw[3][1]),
    .cast_data_o                 (cast_data_pe_2_nw[3][1]),
    .cast_valid_o                (cast_valid_pe_2_nw[3][1]),
    .cast_ready_i                (cast_ready_nw_2_pe[3][1]),
    .merge_data_i                (merge_data_nw_2_pe[3][1]),
    .merge_valid_i               (merge_valid_nw_2_pe[3][1]),
    .merge_ready_o               (merge_ready_pe_2_nw[3][1]),
    .merge_data_o                (merge_data_pe_2_nw[3][1]),
    .merge_valid_o               (merge_valid_pe_2_nw[3][1]),
    .merge_ready_i               (merge_ready_nw_2_pe[3][1])
);


virtual_pe #(
    .isCaster                    (isCaster_3_2)
)vpe_3_2(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[3][2]),
    .cast_valid_i                (cast_valid_nw_2_pe[3][2]),
    .cast_ready_o                (cast_ready_pe_2_nw[3][2]),
    .cast_data_o                 (cast_data_pe_2_nw[3][2]),
    .cast_valid_o                (cast_valid_pe_2_nw[3][2]),
    .cast_ready_i                (cast_ready_nw_2_pe[3][2]),
    .merge_data_i                (merge_data_nw_2_pe[3][2]),
    .merge_valid_i               (merge_valid_nw_2_pe[3][2]),
    .merge_ready_o               (merge_ready_pe_2_nw[3][2]),
    .merge_data_o                (merge_data_pe_2_nw[3][2]),
    .merge_valid_o               (merge_valid_pe_2_nw[3][2]),
    .merge_ready_i               (merge_ready_nw_2_pe[3][2])
);


virtual_pe #(
    .isCaster                    (isCaster_3_3)
)vpe_3_3(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[3][3]),
    .cast_valid_i                (cast_valid_nw_2_pe[3][3]),
    .cast_ready_o                (cast_ready_pe_2_nw[3][3]),
    .cast_data_o                 (cast_data_pe_2_nw[3][3]),
    .cast_valid_o                (cast_valid_pe_2_nw[3][3]),
    .cast_ready_i                (cast_ready_nw_2_pe[3][3]),
    .merge_data_i                (merge_data_nw_2_pe[3][3]),
    .merge_valid_i               (merge_valid_nw_2_pe[3][3]),
    .merge_ready_o               (merge_ready_pe_2_nw[3][3]),
    .merge_data_o                (merge_data_pe_2_nw[3][3]),
    .merge_valid_o               (merge_valid_pe_2_nw[3][3]),
    .merge_ready_i               (merge_ready_nw_2_pe[3][3])
);


virtual_pe #(
    .isCaster                    (isCaster_3_4)
)vpe_3_4(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[3][4]),
    .cast_valid_i                (cast_valid_nw_2_pe[3][4]),
    .cast_ready_o                (cast_ready_pe_2_nw[3][4]),
    .cast_data_o                 (cast_data_pe_2_nw[3][4]),
    .cast_valid_o                (cast_valid_pe_2_nw[3][4]),
    .cast_ready_i                (cast_ready_nw_2_pe[3][4]),
    .merge_data_i                (merge_data_nw_2_pe[3][4]),
    .merge_valid_i               (merge_valid_nw_2_pe[3][4]),
    .merge_ready_o               (merge_ready_pe_2_nw[3][4]),
    .merge_data_o                (merge_data_pe_2_nw[3][4]),
    .merge_valid_o               (merge_valid_pe_2_nw[3][4]),
    .merge_ready_i               (merge_ready_nw_2_pe[3][4])
);


virtual_pe #(
    .isCaster                    (isCaster_3_5)
)vpe_3_5(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[3][5]),
    .cast_valid_i                (cast_valid_nw_2_pe[3][5]),
    .cast_ready_o                (cast_ready_pe_2_nw[3][5]),
    .cast_data_o                 (cast_data_pe_2_nw[3][5]),
    .cast_valid_o                (cast_valid_pe_2_nw[3][5]),
    .cast_ready_i                (cast_ready_nw_2_pe[3][5]),
    .merge_data_i                (merge_data_nw_2_pe[3][5]),
    .merge_valid_i               (merge_valid_nw_2_pe[3][5]),
    .merge_ready_o               (merge_ready_pe_2_nw[3][5]),
    .merge_data_o                (merge_data_pe_2_nw[3][5]),
    .merge_valid_o               (merge_valid_pe_2_nw[3][5]),
    .merge_ready_i               (merge_ready_nw_2_pe[3][5])
);


virtual_pe #(
    .isCaster                    (isCaster_3_6)
)vpe_3_6(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[3][6]),
    .cast_valid_i                (cast_valid_nw_2_pe[3][6]),
    .cast_ready_o                (cast_ready_pe_2_nw[3][6]),
    .cast_data_o                 (cast_data_pe_2_nw[3][6]),
    .cast_valid_o                (cast_valid_pe_2_nw[3][6]),
    .cast_ready_i                (cast_ready_nw_2_pe[3][6]),
    .merge_data_i                (merge_data_nw_2_pe[3][6]),
    .merge_valid_i               (merge_valid_nw_2_pe[3][6]),
    .merge_ready_o               (merge_ready_pe_2_nw[3][6]),
    .merge_data_o                (merge_data_pe_2_nw[3][6]),
    .merge_valid_o               (merge_valid_pe_2_nw[3][6]),
    .merge_ready_i               (merge_ready_nw_2_pe[3][6])
);


virtual_pe #(
    .isCaster                    (isCaster_3_7)
)vpe_3_7(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[3][7]),
    .cast_valid_i                (cast_valid_nw_2_pe[3][7]),
    .cast_ready_o                (cast_ready_pe_2_nw[3][7]),
    .cast_data_o                 (cast_data_pe_2_nw[3][7]),
    .cast_valid_o                (cast_valid_pe_2_nw[3][7]),
    .cast_ready_i                (cast_ready_nw_2_pe[3][7]),
    .merge_data_i                (merge_data_nw_2_pe[3][7]),
    .merge_valid_i               (merge_valid_nw_2_pe[3][7]),
    .merge_ready_o               (merge_ready_pe_2_nw[3][7]),
    .merge_data_o                (merge_data_pe_2_nw[3][7]),
    .merge_valid_o               (merge_valid_pe_2_nw[3][7]),
    .merge_ready_i               (merge_ready_nw_2_pe[3][7])
);


virtual_pe #(
    .isCaster                    (isCaster_4_0)
)vpe_4_0(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[4][0]),
    .cast_valid_i                (cast_valid_nw_2_pe[4][0]),
    .cast_ready_o                (cast_ready_pe_2_nw[4][0]),
    .cast_data_o                 (cast_data_pe_2_nw[4][0]),
    .cast_valid_o                (cast_valid_pe_2_nw[4][0]),
    .cast_ready_i                (cast_ready_nw_2_pe[4][0]),
    .merge_data_i                (merge_data_nw_2_pe[4][0]),
    .merge_valid_i               (merge_valid_nw_2_pe[4][0]),
    .merge_ready_o               (merge_ready_pe_2_nw[4][0]),
    .merge_data_o                (merge_data_pe_2_nw[4][0]),
    .merge_valid_o               (merge_valid_pe_2_nw[4][0]),
    .merge_ready_i               (merge_ready_nw_2_pe[4][0])
);


virtual_pe #(
    .isCaster                    (isCaster_4_1)
)vpe_4_1(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[4][1]),
    .cast_valid_i                (cast_valid_nw_2_pe[4][1]),
    .cast_ready_o                (cast_ready_pe_2_nw[4][1]),
    .cast_data_o                 (cast_data_pe_2_nw[4][1]),
    .cast_valid_o                (cast_valid_pe_2_nw[4][1]),
    .cast_ready_i                (cast_ready_nw_2_pe[4][1]),
    .merge_data_i                (merge_data_nw_2_pe[4][1]),
    .merge_valid_i               (merge_valid_nw_2_pe[4][1]),
    .merge_ready_o               (merge_ready_pe_2_nw[4][1]),
    .merge_data_o                (merge_data_pe_2_nw[4][1]),
    .merge_valid_o               (merge_valid_pe_2_nw[4][1]),
    .merge_ready_i               (merge_ready_nw_2_pe[4][1])
);


virtual_pe #(
    .isCaster                    (isCaster_4_2)
)vpe_4_2(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[4][2]),
    .cast_valid_i                (cast_valid_nw_2_pe[4][2]),
    .cast_ready_o                (cast_ready_pe_2_nw[4][2]),
    .cast_data_o                 (cast_data_pe_2_nw[4][2]),
    .cast_valid_o                (cast_valid_pe_2_nw[4][2]),
    .cast_ready_i                (cast_ready_nw_2_pe[4][2]),
    .merge_data_i                (merge_data_nw_2_pe[4][2]),
    .merge_valid_i               (merge_valid_nw_2_pe[4][2]),
    .merge_ready_o               (merge_ready_pe_2_nw[4][2]),
    .merge_data_o                (merge_data_pe_2_nw[4][2]),
    .merge_valid_o               (merge_valid_pe_2_nw[4][2]),
    .merge_ready_i               (merge_ready_nw_2_pe[4][2])
);


virtual_pe #(
    .isCaster                    (isCaster_4_3)
)vpe_4_3(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[4][3]),
    .cast_valid_i                (cast_valid_nw_2_pe[4][3]),
    .cast_ready_o                (cast_ready_pe_2_nw[4][3]),
    .cast_data_o                 (cast_data_pe_2_nw[4][3]),
    .cast_valid_o                (cast_valid_pe_2_nw[4][3]),
    .cast_ready_i                (cast_ready_nw_2_pe[4][3]),
    .merge_data_i                (merge_data_nw_2_pe[4][3]),
    .merge_valid_i               (merge_valid_nw_2_pe[4][3]),
    .merge_ready_o               (merge_ready_pe_2_nw[4][3]),
    .merge_data_o                (merge_data_pe_2_nw[4][3]),
    .merge_valid_o               (merge_valid_pe_2_nw[4][3]),
    .merge_ready_i               (merge_ready_nw_2_pe[4][3])
);


virtual_pe #(
    .isCaster                    (isCaster_4_4)
)vpe_4_4(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[4][4]),
    .cast_valid_i                (cast_valid_nw_2_pe[4][4]),
    .cast_ready_o                (cast_ready_pe_2_nw[4][4]),
    .cast_data_o                 (cast_data_pe_2_nw[4][4]),
    .cast_valid_o                (cast_valid_pe_2_nw[4][4]),
    .cast_ready_i                (cast_ready_nw_2_pe[4][4]),
    .merge_data_i                (merge_data_nw_2_pe[4][4]),
    .merge_valid_i               (merge_valid_nw_2_pe[4][4]),
    .merge_ready_o               (merge_ready_pe_2_nw[4][4]),
    .merge_data_o                (merge_data_pe_2_nw[4][4]),
    .merge_valid_o               (merge_valid_pe_2_nw[4][4]),
    .merge_ready_i               (merge_ready_nw_2_pe[4][4])
);


virtual_pe #(
    .isCaster                    (isCaster_4_5)
)vpe_4_5(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[4][5]),
    .cast_valid_i                (cast_valid_nw_2_pe[4][5]),
    .cast_ready_o                (cast_ready_pe_2_nw[4][5]),
    .cast_data_o                 (cast_data_pe_2_nw[4][5]),
    .cast_valid_o                (cast_valid_pe_2_nw[4][5]),
    .cast_ready_i                (cast_ready_nw_2_pe[4][5]),
    .merge_data_i                (merge_data_nw_2_pe[4][5]),
    .merge_valid_i               (merge_valid_nw_2_pe[4][5]),
    .merge_ready_o               (merge_ready_pe_2_nw[4][5]),
    .merge_data_o                (merge_data_pe_2_nw[4][5]),
    .merge_valid_o               (merge_valid_pe_2_nw[4][5]),
    .merge_ready_i               (merge_ready_nw_2_pe[4][5])
);


virtual_pe #(
    .isCaster                    (isCaster_4_6)
)vpe_4_6(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[4][6]),
    .cast_valid_i                (cast_valid_nw_2_pe[4][6]),
    .cast_ready_o                (cast_ready_pe_2_nw[4][6]),
    .cast_data_o                 (cast_data_pe_2_nw[4][6]),
    .cast_valid_o                (cast_valid_pe_2_nw[4][6]),
    .cast_ready_i                (cast_ready_nw_2_pe[4][6]),
    .merge_data_i                (merge_data_nw_2_pe[4][6]),
    .merge_valid_i               (merge_valid_nw_2_pe[4][6]),
    .merge_ready_o               (merge_ready_pe_2_nw[4][6]),
    .merge_data_o                (merge_data_pe_2_nw[4][6]),
    .merge_valid_o               (merge_valid_pe_2_nw[4][6]),
    .merge_ready_i               (merge_ready_nw_2_pe[4][6])
);


virtual_pe #(
    .isCaster                    (isCaster_4_7)
)vpe_4_7(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[4][7]),
    .cast_valid_i                (cast_valid_nw_2_pe[4][7]),
    .cast_ready_o                (cast_ready_pe_2_nw[4][7]),
    .cast_data_o                 (cast_data_pe_2_nw[4][7]),
    .cast_valid_o                (cast_valid_pe_2_nw[4][7]),
    .cast_ready_i                (cast_ready_nw_2_pe[4][7]),
    .merge_data_i                (merge_data_nw_2_pe[4][7]),
    .merge_valid_i               (merge_valid_nw_2_pe[4][7]),
    .merge_ready_o               (merge_ready_pe_2_nw[4][7]),
    .merge_data_o                (merge_data_pe_2_nw[4][7]),
    .merge_valid_o               (merge_valid_pe_2_nw[4][7]),
    .merge_ready_i               (merge_ready_nw_2_pe[4][7])
);


virtual_pe #(
    .isCaster                    (isCaster_5_0)
)vpe_5_0(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[5][0]),
    .cast_valid_i                (cast_valid_nw_2_pe[5][0]),
    .cast_ready_o                (cast_ready_pe_2_nw[5][0]),
    .cast_data_o                 (cast_data_pe_2_nw[5][0]),
    .cast_valid_o                (cast_valid_pe_2_nw[5][0]),
    .cast_ready_i                (cast_ready_nw_2_pe[5][0]),
    .merge_data_i                (merge_data_nw_2_pe[5][0]),
    .merge_valid_i               (merge_valid_nw_2_pe[5][0]),
    .merge_ready_o               (merge_ready_pe_2_nw[5][0]),
    .merge_data_o                (merge_data_pe_2_nw[5][0]),
    .merge_valid_o               (merge_valid_pe_2_nw[5][0]),
    .merge_ready_i               (merge_ready_nw_2_pe[5][0])
);


virtual_pe #(
    .isCaster                    (isCaster_5_1)
)vpe_5_1(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[5][1]),
    .cast_valid_i                (cast_valid_nw_2_pe[5][1]),
    .cast_ready_o                (cast_ready_pe_2_nw[5][1]),
    .cast_data_o                 (cast_data_pe_2_nw[5][1]),
    .cast_valid_o                (cast_valid_pe_2_nw[5][1]),
    .cast_ready_i                (cast_ready_nw_2_pe[5][1]),
    .merge_data_i                (merge_data_nw_2_pe[5][1]),
    .merge_valid_i               (merge_valid_nw_2_pe[5][1]),
    .merge_ready_o               (merge_ready_pe_2_nw[5][1]),
    .merge_data_o                (merge_data_pe_2_nw[5][1]),
    .merge_valid_o               (merge_valid_pe_2_nw[5][1]),
    .merge_ready_i               (merge_ready_nw_2_pe[5][1])
);


virtual_pe #(
    .isCaster                    (isCaster_5_2)
)vpe_5_2(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[5][2]),
    .cast_valid_i                (cast_valid_nw_2_pe[5][2]),
    .cast_ready_o                (cast_ready_pe_2_nw[5][2]),
    .cast_data_o                 (cast_data_pe_2_nw[5][2]),
    .cast_valid_o                (cast_valid_pe_2_nw[5][2]),
    .cast_ready_i                (cast_ready_nw_2_pe[5][2]),
    .merge_data_i                (merge_data_nw_2_pe[5][2]),
    .merge_valid_i               (merge_valid_nw_2_pe[5][2]),
    .merge_ready_o               (merge_ready_pe_2_nw[5][2]),
    .merge_data_o                (merge_data_pe_2_nw[5][2]),
    .merge_valid_o               (merge_valid_pe_2_nw[5][2]),
    .merge_ready_i               (merge_ready_nw_2_pe[5][2])
);


virtual_pe #(
    .isCaster                    (isCaster_5_3)
)vpe_5_3(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[5][3]),
    .cast_valid_i                (cast_valid_nw_2_pe[5][3]),
    .cast_ready_o                (cast_ready_pe_2_nw[5][3]),
    .cast_data_o                 (cast_data_pe_2_nw[5][3]),
    .cast_valid_o                (cast_valid_pe_2_nw[5][3]),
    .cast_ready_i                (cast_ready_nw_2_pe[5][3]),
    .merge_data_i                (merge_data_nw_2_pe[5][3]),
    .merge_valid_i               (merge_valid_nw_2_pe[5][3]),
    .merge_ready_o               (merge_ready_pe_2_nw[5][3]),
    .merge_data_o                (merge_data_pe_2_nw[5][3]),
    .merge_valid_o               (merge_valid_pe_2_nw[5][3]),
    .merge_ready_i               (merge_ready_nw_2_pe[5][3])
);


virtual_pe #(
    .isCaster                    (isCaster_5_4)
)vpe_5_4(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[5][4]),
    .cast_valid_i                (cast_valid_nw_2_pe[5][4]),
    .cast_ready_o                (cast_ready_pe_2_nw[5][4]),
    .cast_data_o                 (cast_data_pe_2_nw[5][4]),
    .cast_valid_o                (cast_valid_pe_2_nw[5][4]),
    .cast_ready_i                (cast_ready_nw_2_pe[5][4]),
    .merge_data_i                (merge_data_nw_2_pe[5][4]),
    .merge_valid_i               (merge_valid_nw_2_pe[5][4]),
    .merge_ready_o               (merge_ready_pe_2_nw[5][4]),
    .merge_data_o                (merge_data_pe_2_nw[5][4]),
    .merge_valid_o               (merge_valid_pe_2_nw[5][4]),
    .merge_ready_i               (merge_ready_nw_2_pe[5][4])
);


virtual_pe #(
    .isCaster                    (isCaster_5_5)
)vpe_5_5(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[5][5]),
    .cast_valid_i                (cast_valid_nw_2_pe[5][5]),
    .cast_ready_o                (cast_ready_pe_2_nw[5][5]),
    .cast_data_o                 (cast_data_pe_2_nw[5][5]),
    .cast_valid_o                (cast_valid_pe_2_nw[5][5]),
    .cast_ready_i                (cast_ready_nw_2_pe[5][5]),
    .merge_data_i                (merge_data_nw_2_pe[5][5]),
    .merge_valid_i               (merge_valid_nw_2_pe[5][5]),
    .merge_ready_o               (merge_ready_pe_2_nw[5][5]),
    .merge_data_o                (merge_data_pe_2_nw[5][5]),
    .merge_valid_o               (merge_valid_pe_2_nw[5][5]),
    .merge_ready_i               (merge_ready_nw_2_pe[5][5])
);


virtual_pe #(
    .isCaster                    (isCaster_5_6)
)vpe_5_6(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[5][6]),
    .cast_valid_i                (cast_valid_nw_2_pe[5][6]),
    .cast_ready_o                (cast_ready_pe_2_nw[5][6]),
    .cast_data_o                 (cast_data_pe_2_nw[5][6]),
    .cast_valid_o                (cast_valid_pe_2_nw[5][6]),
    .cast_ready_i                (cast_ready_nw_2_pe[5][6]),
    .merge_data_i                (merge_data_nw_2_pe[5][6]),
    .merge_valid_i               (merge_valid_nw_2_pe[5][6]),
    .merge_ready_o               (merge_ready_pe_2_nw[5][6]),
    .merge_data_o                (merge_data_pe_2_nw[5][6]),
    .merge_valid_o               (merge_valid_pe_2_nw[5][6]),
    .merge_ready_i               (merge_ready_nw_2_pe[5][6])
);


virtual_pe #(
    .isCaster                    (isCaster_5_7)
)vpe_5_7(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[5][7]),
    .cast_valid_i                (cast_valid_nw_2_pe[5][7]),
    .cast_ready_o                (cast_ready_pe_2_nw[5][7]),
    .cast_data_o                 (cast_data_pe_2_nw[5][7]),
    .cast_valid_o                (cast_valid_pe_2_nw[5][7]),
    .cast_ready_i                (cast_ready_nw_2_pe[5][7]),
    .merge_data_i                (merge_data_nw_2_pe[5][7]),
    .merge_valid_i               (merge_valid_nw_2_pe[5][7]),
    .merge_ready_o               (merge_ready_pe_2_nw[5][7]),
    .merge_data_o                (merge_data_pe_2_nw[5][7]),
    .merge_valid_o               (merge_valid_pe_2_nw[5][7]),
    .merge_ready_i               (merge_ready_nw_2_pe[5][7])
);


virtual_pe #(
    .isCaster                    (isCaster_6_0)
)vpe_6_0(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[6][0]),
    .cast_valid_i                (cast_valid_nw_2_pe[6][0]),
    .cast_ready_o                (cast_ready_pe_2_nw[6][0]),
    .cast_data_o                 (cast_data_pe_2_nw[6][0]),
    .cast_valid_o                (cast_valid_pe_2_nw[6][0]),
    .cast_ready_i                (cast_ready_nw_2_pe[6][0]),
    .merge_data_i                (merge_data_nw_2_pe[6][0]),
    .merge_valid_i               (merge_valid_nw_2_pe[6][0]),
    .merge_ready_o               (merge_ready_pe_2_nw[6][0]),
    .merge_data_o                (merge_data_pe_2_nw[6][0]),
    .merge_valid_o               (merge_valid_pe_2_nw[6][0]),
    .merge_ready_i               (merge_ready_nw_2_pe[6][0])
);


virtual_pe #(
    .isCaster                    (isCaster_6_1)
)vpe_6_1(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[6][1]),
    .cast_valid_i                (cast_valid_nw_2_pe[6][1]),
    .cast_ready_o                (cast_ready_pe_2_nw[6][1]),
    .cast_data_o                 (cast_data_pe_2_nw[6][1]),
    .cast_valid_o                (cast_valid_pe_2_nw[6][1]),
    .cast_ready_i                (cast_ready_nw_2_pe[6][1]),
    .merge_data_i                (merge_data_nw_2_pe[6][1]),
    .merge_valid_i               (merge_valid_nw_2_pe[6][1]),
    .merge_ready_o               (merge_ready_pe_2_nw[6][1]),
    .merge_data_o                (merge_data_pe_2_nw[6][1]),
    .merge_valid_o               (merge_valid_pe_2_nw[6][1]),
    .merge_ready_i               (merge_ready_nw_2_pe[6][1])
);


virtual_pe #(
    .isCaster                    (isCaster_6_2)
)vpe_6_2(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[6][2]),
    .cast_valid_i                (cast_valid_nw_2_pe[6][2]),
    .cast_ready_o                (cast_ready_pe_2_nw[6][2]),
    .cast_data_o                 (cast_data_pe_2_nw[6][2]),
    .cast_valid_o                (cast_valid_pe_2_nw[6][2]),
    .cast_ready_i                (cast_ready_nw_2_pe[6][2]),
    .merge_data_i                (merge_data_nw_2_pe[6][2]),
    .merge_valid_i               (merge_valid_nw_2_pe[6][2]),
    .merge_ready_o               (merge_ready_pe_2_nw[6][2]),
    .merge_data_o                (merge_data_pe_2_nw[6][2]),
    .merge_valid_o               (merge_valid_pe_2_nw[6][2]),
    .merge_ready_i               (merge_ready_nw_2_pe[6][2])
);


virtual_pe #(
    .isCaster                    (isCaster_6_3)
)vpe_6_3(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[6][3]),
    .cast_valid_i                (cast_valid_nw_2_pe[6][3]),
    .cast_ready_o                (cast_ready_pe_2_nw[6][3]),
    .cast_data_o                 (cast_data_pe_2_nw[6][3]),
    .cast_valid_o                (cast_valid_pe_2_nw[6][3]),
    .cast_ready_i                (cast_ready_nw_2_pe[6][3]),
    .merge_data_i                (merge_data_nw_2_pe[6][3]),
    .merge_valid_i               (merge_valid_nw_2_pe[6][3]),
    .merge_ready_o               (merge_ready_pe_2_nw[6][3]),
    .merge_data_o                (merge_data_pe_2_nw[6][3]),
    .merge_valid_o               (merge_valid_pe_2_nw[6][3]),
    .merge_ready_i               (merge_ready_nw_2_pe[6][3])
);


virtual_pe #(
    .isCaster                    (isCaster_6_4)
)vpe_6_4(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[6][4]),
    .cast_valid_i                (cast_valid_nw_2_pe[6][4]),
    .cast_ready_o                (cast_ready_pe_2_nw[6][4]),
    .cast_data_o                 (cast_data_pe_2_nw[6][4]),
    .cast_valid_o                (cast_valid_pe_2_nw[6][4]),
    .cast_ready_i                (cast_ready_nw_2_pe[6][4]),
    .merge_data_i                (merge_data_nw_2_pe[6][4]),
    .merge_valid_i               (merge_valid_nw_2_pe[6][4]),
    .merge_ready_o               (merge_ready_pe_2_nw[6][4]),
    .merge_data_o                (merge_data_pe_2_nw[6][4]),
    .merge_valid_o               (merge_valid_pe_2_nw[6][4]),
    .merge_ready_i               (merge_ready_nw_2_pe[6][4])
);


virtual_pe #(
    .isCaster                    (isCaster_6_5)
)vpe_6_5(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[6][5]),
    .cast_valid_i                (cast_valid_nw_2_pe[6][5]),
    .cast_ready_o                (cast_ready_pe_2_nw[6][5]),
    .cast_data_o                 (cast_data_pe_2_nw[6][5]),
    .cast_valid_o                (cast_valid_pe_2_nw[6][5]),
    .cast_ready_i                (cast_ready_nw_2_pe[6][5]),
    .merge_data_i                (merge_data_nw_2_pe[6][5]),
    .merge_valid_i               (merge_valid_nw_2_pe[6][5]),
    .merge_ready_o               (merge_ready_pe_2_nw[6][5]),
    .merge_data_o                (merge_data_pe_2_nw[6][5]),
    .merge_valid_o               (merge_valid_pe_2_nw[6][5]),
    .merge_ready_i               (merge_ready_nw_2_pe[6][5])
);


virtual_pe #(
    .isCaster                    (isCaster_6_6)
)vpe_6_6(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[6][6]),
    .cast_valid_i                (cast_valid_nw_2_pe[6][6]),
    .cast_ready_o                (cast_ready_pe_2_nw[6][6]),
    .cast_data_o                 (cast_data_pe_2_nw[6][6]),
    .cast_valid_o                (cast_valid_pe_2_nw[6][6]),
    .cast_ready_i                (cast_ready_nw_2_pe[6][6]),
    .merge_data_i                (merge_data_nw_2_pe[6][6]),
    .merge_valid_i               (merge_valid_nw_2_pe[6][6]),
    .merge_ready_o               (merge_ready_pe_2_nw[6][6]),
    .merge_data_o                (merge_data_pe_2_nw[6][6]),
    .merge_valid_o               (merge_valid_pe_2_nw[6][6]),
    .merge_ready_i               (merge_ready_nw_2_pe[6][6])
);


virtual_pe #(
    .isCaster                    (isCaster_6_7)
)vpe_6_7(
    .clk                         (clk),
    .rstn                        (rstn),
    .cast_data_i                 (cast_data_nw_2_pe[6][7]),
    .cast_valid_i                (cast_valid_nw_2_pe[6][7]),
    .cast_ready_o                (cast_ready_pe_2_nw[6][7]),
    .cast_data_o                 (cast_data_pe_2_nw[6][7]),
    .cast_valid_o                (cast_valid_pe_2_nw[6][7]),
    .cast_ready_i                (cast_ready_nw_2_pe[6][7]),
    .merge_data_i                (merge_data_nw_2_pe[6][7]),
    .merge_valid_i               (merge_valid_nw_2_pe[6][7]),
    .merge_ready_o               (merge_ready_pe_2_nw[6][7]),
    .merge_data_o                (merge_data_pe_2_nw[6][7]),
    .merge_valid_o               (merge_valid_pe_2_nw[6][7]),
    .merge_ready_i               (merge_ready_nw_2_pe[6][7])
);

endmodule
