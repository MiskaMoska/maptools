
//Merge Network
//Width: 10
//Height:25
`include "params.svh"
`include "merge_network_config.svh"

module merge_network(
    input       wire                            clk,
    input       wire                            rstn,

    //router local ports
    input       wire        [`DW-1:0]           data_i[`NOC_WIDTH][`NOC_HEIGHT],
    input       wire                            valid_i[`NOC_WIDTH][`NOC_HEIGHT],
    output      reg                             ready_o[`NOC_WIDTH][`NOC_HEIGHT],

    output      reg         [`DW-1:0]           data_o[`NOC_WIDTH][`NOC_HEIGHT],
    output      reg                             valid_o[`NOC_WIDTH][`NOC_HEIGHT],
    input       wire                            ready_i[`NOC_WIDTH][`NOC_HEIGHT]
);

reg [`DW-1:0] data_i_0_0[5];
reg valid_i_0_0[5], ready_i_0_0[5];    
wire [`DW-1:0] data_o_0_0[5];
wire valid_o_0_0[5], ready_o_0_0[5];        

reg [`DW-1:0] data_i_0_1[5];
reg valid_i_0_1[5], ready_i_0_1[5];    
wire [`DW-1:0] data_o_0_1[5];
wire valid_o_0_1[5], ready_o_0_1[5];        

reg [`DW-1:0] data_i_0_2[5];
reg valid_i_0_2[5], ready_i_0_2[5];    
wire [`DW-1:0] data_o_0_2[5];
wire valid_o_0_2[5], ready_o_0_2[5];        

reg [`DW-1:0] data_i_0_3[5];
reg valid_i_0_3[5], ready_i_0_3[5];    
wire [`DW-1:0] data_o_0_3[5];
wire valid_o_0_3[5], ready_o_0_3[5];        

reg [`DW-1:0] data_i_0_4[5];
reg valid_i_0_4[5], ready_i_0_4[5];    
wire [`DW-1:0] data_o_0_4[5];
wire valid_o_0_4[5], ready_o_0_4[5];        

reg [`DW-1:0] data_i_0_5[5];
reg valid_i_0_5[5], ready_i_0_5[5];    
wire [`DW-1:0] data_o_0_5[5];
wire valid_o_0_5[5], ready_o_0_5[5];        

reg [`DW-1:0] data_i_0_6[5];
reg valid_i_0_6[5], ready_i_0_6[5];    
wire [`DW-1:0] data_o_0_6[5];
wire valid_o_0_6[5], ready_o_0_6[5];        

reg [`DW-1:0] data_i_0_7[5];
reg valid_i_0_7[5], ready_i_0_7[5];    
wire [`DW-1:0] data_o_0_7[5];
wire valid_o_0_7[5], ready_o_0_7[5];        

reg [`DW-1:0] data_i_0_8[5];
reg valid_i_0_8[5], ready_i_0_8[5];    
wire [`DW-1:0] data_o_0_8[5];
wire valid_o_0_8[5], ready_o_0_8[5];        

reg [`DW-1:0] data_i_0_9[5];
reg valid_i_0_9[5], ready_i_0_9[5];    
wire [`DW-1:0] data_o_0_9[5];
wire valid_o_0_9[5], ready_o_0_9[5];        

reg [`DW-1:0] data_i_0_10[5];
reg valid_i_0_10[5], ready_i_0_10[5];    
wire [`DW-1:0] data_o_0_10[5];
wire valid_o_0_10[5], ready_o_0_10[5];        

reg [`DW-1:0] data_i_0_11[5];
reg valid_i_0_11[5], ready_i_0_11[5];    
wire [`DW-1:0] data_o_0_11[5];
wire valid_o_0_11[5], ready_o_0_11[5];        

reg [`DW-1:0] data_i_0_12[5];
reg valid_i_0_12[5], ready_i_0_12[5];    
wire [`DW-1:0] data_o_0_12[5];
wire valid_o_0_12[5], ready_o_0_12[5];        

reg [`DW-1:0] data_i_0_13[5];
reg valid_i_0_13[5], ready_i_0_13[5];    
wire [`DW-1:0] data_o_0_13[5];
wire valid_o_0_13[5], ready_o_0_13[5];        

reg [`DW-1:0] data_i_0_14[5];
reg valid_i_0_14[5], ready_i_0_14[5];    
wire [`DW-1:0] data_o_0_14[5];
wire valid_o_0_14[5], ready_o_0_14[5];        

reg [`DW-1:0] data_i_0_15[5];
reg valid_i_0_15[5], ready_i_0_15[5];    
wire [`DW-1:0] data_o_0_15[5];
wire valid_o_0_15[5], ready_o_0_15[5];        

reg [`DW-1:0] data_i_0_16[5];
reg valid_i_0_16[5], ready_i_0_16[5];    
wire [`DW-1:0] data_o_0_16[5];
wire valid_o_0_16[5], ready_o_0_16[5];        

reg [`DW-1:0] data_i_0_17[5];
reg valid_i_0_17[5], ready_i_0_17[5];    
wire [`DW-1:0] data_o_0_17[5];
wire valid_o_0_17[5], ready_o_0_17[5];        

reg [`DW-1:0] data_i_0_18[5];
reg valid_i_0_18[5], ready_i_0_18[5];    
wire [`DW-1:0] data_o_0_18[5];
wire valid_o_0_18[5], ready_o_0_18[5];        

reg [`DW-1:0] data_i_0_19[5];
reg valid_i_0_19[5], ready_i_0_19[5];    
wire [`DW-1:0] data_o_0_19[5];
wire valid_o_0_19[5], ready_o_0_19[5];        

reg [`DW-1:0] data_i_0_20[5];
reg valid_i_0_20[5], ready_i_0_20[5];    
wire [`DW-1:0] data_o_0_20[5];
wire valid_o_0_20[5], ready_o_0_20[5];        

reg [`DW-1:0] data_i_0_21[5];
reg valid_i_0_21[5], ready_i_0_21[5];    
wire [`DW-1:0] data_o_0_21[5];
wire valid_o_0_21[5], ready_o_0_21[5];        

reg [`DW-1:0] data_i_0_22[5];
reg valid_i_0_22[5], ready_i_0_22[5];    
wire [`DW-1:0] data_o_0_22[5];
wire valid_o_0_22[5], ready_o_0_22[5];        

reg [`DW-1:0] data_i_0_23[5];
reg valid_i_0_23[5], ready_i_0_23[5];    
wire [`DW-1:0] data_o_0_23[5];
wire valid_o_0_23[5], ready_o_0_23[5];        

reg [`DW-1:0] data_i_0_24[5];
reg valid_i_0_24[5], ready_i_0_24[5];    
wire [`DW-1:0] data_o_0_24[5];
wire valid_o_0_24[5], ready_o_0_24[5];        

reg [`DW-1:0] data_i_1_0[5];
reg valid_i_1_0[5], ready_i_1_0[5];    
wire [`DW-1:0] data_o_1_0[5];
wire valid_o_1_0[5], ready_o_1_0[5];        

reg [`DW-1:0] data_i_1_1[5];
reg valid_i_1_1[5], ready_i_1_1[5];    
wire [`DW-1:0] data_o_1_1[5];
wire valid_o_1_1[5], ready_o_1_1[5];        

reg [`DW-1:0] data_i_1_2[5];
reg valid_i_1_2[5], ready_i_1_2[5];    
wire [`DW-1:0] data_o_1_2[5];
wire valid_o_1_2[5], ready_o_1_2[5];        

reg [`DW-1:0] data_i_1_3[5];
reg valid_i_1_3[5], ready_i_1_3[5];    
wire [`DW-1:0] data_o_1_3[5];
wire valid_o_1_3[5], ready_o_1_3[5];        

reg [`DW-1:0] data_i_1_4[5];
reg valid_i_1_4[5], ready_i_1_4[5];    
wire [`DW-1:0] data_o_1_4[5];
wire valid_o_1_4[5], ready_o_1_4[5];        

reg [`DW-1:0] data_i_1_5[5];
reg valid_i_1_5[5], ready_i_1_5[5];    
wire [`DW-1:0] data_o_1_5[5];
wire valid_o_1_5[5], ready_o_1_5[5];        

reg [`DW-1:0] data_i_1_6[5];
reg valid_i_1_6[5], ready_i_1_6[5];    
wire [`DW-1:0] data_o_1_6[5];
wire valid_o_1_6[5], ready_o_1_6[5];        

reg [`DW-1:0] data_i_1_7[5];
reg valid_i_1_7[5], ready_i_1_7[5];    
wire [`DW-1:0] data_o_1_7[5];
wire valid_o_1_7[5], ready_o_1_7[5];        

reg [`DW-1:0] data_i_1_8[5];
reg valid_i_1_8[5], ready_i_1_8[5];    
wire [`DW-1:0] data_o_1_8[5];
wire valid_o_1_8[5], ready_o_1_8[5];        

reg [`DW-1:0] data_i_1_9[5];
reg valid_i_1_9[5], ready_i_1_9[5];    
wire [`DW-1:0] data_o_1_9[5];
wire valid_o_1_9[5], ready_o_1_9[5];        

reg [`DW-1:0] data_i_1_10[5];
reg valid_i_1_10[5], ready_i_1_10[5];    
wire [`DW-1:0] data_o_1_10[5];
wire valid_o_1_10[5], ready_o_1_10[5];        

reg [`DW-1:0] data_i_1_11[5];
reg valid_i_1_11[5], ready_i_1_11[5];    
wire [`DW-1:0] data_o_1_11[5];
wire valid_o_1_11[5], ready_o_1_11[5];        

reg [`DW-1:0] data_i_1_12[5];
reg valid_i_1_12[5], ready_i_1_12[5];    
wire [`DW-1:0] data_o_1_12[5];
wire valid_o_1_12[5], ready_o_1_12[5];        

reg [`DW-1:0] data_i_1_13[5];
reg valid_i_1_13[5], ready_i_1_13[5];    
wire [`DW-1:0] data_o_1_13[5];
wire valid_o_1_13[5], ready_o_1_13[5];        

reg [`DW-1:0] data_i_1_14[5];
reg valid_i_1_14[5], ready_i_1_14[5];    
wire [`DW-1:0] data_o_1_14[5];
wire valid_o_1_14[5], ready_o_1_14[5];        

reg [`DW-1:0] data_i_1_15[5];
reg valid_i_1_15[5], ready_i_1_15[5];    
wire [`DW-1:0] data_o_1_15[5];
wire valid_o_1_15[5], ready_o_1_15[5];        

reg [`DW-1:0] data_i_1_16[5];
reg valid_i_1_16[5], ready_i_1_16[5];    
wire [`DW-1:0] data_o_1_16[5];
wire valid_o_1_16[5], ready_o_1_16[5];        

reg [`DW-1:0] data_i_1_17[5];
reg valid_i_1_17[5], ready_i_1_17[5];    
wire [`DW-1:0] data_o_1_17[5];
wire valid_o_1_17[5], ready_o_1_17[5];        

reg [`DW-1:0] data_i_1_18[5];
reg valid_i_1_18[5], ready_i_1_18[5];    
wire [`DW-1:0] data_o_1_18[5];
wire valid_o_1_18[5], ready_o_1_18[5];        

reg [`DW-1:0] data_i_1_19[5];
reg valid_i_1_19[5], ready_i_1_19[5];    
wire [`DW-1:0] data_o_1_19[5];
wire valid_o_1_19[5], ready_o_1_19[5];        

reg [`DW-1:0] data_i_1_20[5];
reg valid_i_1_20[5], ready_i_1_20[5];    
wire [`DW-1:0] data_o_1_20[5];
wire valid_o_1_20[5], ready_o_1_20[5];        

reg [`DW-1:0] data_i_1_21[5];
reg valid_i_1_21[5], ready_i_1_21[5];    
wire [`DW-1:0] data_o_1_21[5];
wire valid_o_1_21[5], ready_o_1_21[5];        

reg [`DW-1:0] data_i_1_22[5];
reg valid_i_1_22[5], ready_i_1_22[5];    
wire [`DW-1:0] data_o_1_22[5];
wire valid_o_1_22[5], ready_o_1_22[5];        

reg [`DW-1:0] data_i_1_23[5];
reg valid_i_1_23[5], ready_i_1_23[5];    
wire [`DW-1:0] data_o_1_23[5];
wire valid_o_1_23[5], ready_o_1_23[5];        

reg [`DW-1:0] data_i_1_24[5];
reg valid_i_1_24[5], ready_i_1_24[5];    
wire [`DW-1:0] data_o_1_24[5];
wire valid_o_1_24[5], ready_o_1_24[5];        

reg [`DW-1:0] data_i_2_0[5];
reg valid_i_2_0[5], ready_i_2_0[5];    
wire [`DW-1:0] data_o_2_0[5];
wire valid_o_2_0[5], ready_o_2_0[5];        

reg [`DW-1:0] data_i_2_1[5];
reg valid_i_2_1[5], ready_i_2_1[5];    
wire [`DW-1:0] data_o_2_1[5];
wire valid_o_2_1[5], ready_o_2_1[5];        

reg [`DW-1:0] data_i_2_2[5];
reg valid_i_2_2[5], ready_i_2_2[5];    
wire [`DW-1:0] data_o_2_2[5];
wire valid_o_2_2[5], ready_o_2_2[5];        

reg [`DW-1:0] data_i_2_3[5];
reg valid_i_2_3[5], ready_i_2_3[5];    
wire [`DW-1:0] data_o_2_3[5];
wire valid_o_2_3[5], ready_o_2_3[5];        

reg [`DW-1:0] data_i_2_4[5];
reg valid_i_2_4[5], ready_i_2_4[5];    
wire [`DW-1:0] data_o_2_4[5];
wire valid_o_2_4[5], ready_o_2_4[5];        

reg [`DW-1:0] data_i_2_5[5];
reg valid_i_2_5[5], ready_i_2_5[5];    
wire [`DW-1:0] data_o_2_5[5];
wire valid_o_2_5[5], ready_o_2_5[5];        

reg [`DW-1:0] data_i_2_6[5];
reg valid_i_2_6[5], ready_i_2_6[5];    
wire [`DW-1:0] data_o_2_6[5];
wire valid_o_2_6[5], ready_o_2_6[5];        

reg [`DW-1:0] data_i_2_7[5];
reg valid_i_2_7[5], ready_i_2_7[5];    
wire [`DW-1:0] data_o_2_7[5];
wire valid_o_2_7[5], ready_o_2_7[5];        

reg [`DW-1:0] data_i_2_8[5];
reg valid_i_2_8[5], ready_i_2_8[5];    
wire [`DW-1:0] data_o_2_8[5];
wire valid_o_2_8[5], ready_o_2_8[5];        

reg [`DW-1:0] data_i_2_9[5];
reg valid_i_2_9[5], ready_i_2_9[5];    
wire [`DW-1:0] data_o_2_9[5];
wire valid_o_2_9[5], ready_o_2_9[5];        

reg [`DW-1:0] data_i_2_10[5];
reg valid_i_2_10[5], ready_i_2_10[5];    
wire [`DW-1:0] data_o_2_10[5];
wire valid_o_2_10[5], ready_o_2_10[5];        

reg [`DW-1:0] data_i_2_11[5];
reg valid_i_2_11[5], ready_i_2_11[5];    
wire [`DW-1:0] data_o_2_11[5];
wire valid_o_2_11[5], ready_o_2_11[5];        

reg [`DW-1:0] data_i_2_12[5];
reg valid_i_2_12[5], ready_i_2_12[5];    
wire [`DW-1:0] data_o_2_12[5];
wire valid_o_2_12[5], ready_o_2_12[5];        

reg [`DW-1:0] data_i_2_13[5];
reg valid_i_2_13[5], ready_i_2_13[5];    
wire [`DW-1:0] data_o_2_13[5];
wire valid_o_2_13[5], ready_o_2_13[5];        

reg [`DW-1:0] data_i_2_14[5];
reg valid_i_2_14[5], ready_i_2_14[5];    
wire [`DW-1:0] data_o_2_14[5];
wire valid_o_2_14[5], ready_o_2_14[5];        

reg [`DW-1:0] data_i_2_15[5];
reg valid_i_2_15[5], ready_i_2_15[5];    
wire [`DW-1:0] data_o_2_15[5];
wire valid_o_2_15[5], ready_o_2_15[5];        

reg [`DW-1:0] data_i_2_16[5];
reg valid_i_2_16[5], ready_i_2_16[5];    
wire [`DW-1:0] data_o_2_16[5];
wire valid_o_2_16[5], ready_o_2_16[5];        

reg [`DW-1:0] data_i_2_17[5];
reg valid_i_2_17[5], ready_i_2_17[5];    
wire [`DW-1:0] data_o_2_17[5];
wire valid_o_2_17[5], ready_o_2_17[5];        

reg [`DW-1:0] data_i_2_18[5];
reg valid_i_2_18[5], ready_i_2_18[5];    
wire [`DW-1:0] data_o_2_18[5];
wire valid_o_2_18[5], ready_o_2_18[5];        

reg [`DW-1:0] data_i_2_19[5];
reg valid_i_2_19[5], ready_i_2_19[5];    
wire [`DW-1:0] data_o_2_19[5];
wire valid_o_2_19[5], ready_o_2_19[5];        

reg [`DW-1:0] data_i_2_20[5];
reg valid_i_2_20[5], ready_i_2_20[5];    
wire [`DW-1:0] data_o_2_20[5];
wire valid_o_2_20[5], ready_o_2_20[5];        

reg [`DW-1:0] data_i_2_21[5];
reg valid_i_2_21[5], ready_i_2_21[5];    
wire [`DW-1:0] data_o_2_21[5];
wire valid_o_2_21[5], ready_o_2_21[5];        

reg [`DW-1:0] data_i_2_22[5];
reg valid_i_2_22[5], ready_i_2_22[5];    
wire [`DW-1:0] data_o_2_22[5];
wire valid_o_2_22[5], ready_o_2_22[5];        

reg [`DW-1:0] data_i_2_23[5];
reg valid_i_2_23[5], ready_i_2_23[5];    
wire [`DW-1:0] data_o_2_23[5];
wire valid_o_2_23[5], ready_o_2_23[5];        

reg [`DW-1:0] data_i_2_24[5];
reg valid_i_2_24[5], ready_i_2_24[5];    
wire [`DW-1:0] data_o_2_24[5];
wire valid_o_2_24[5], ready_o_2_24[5];        

reg [`DW-1:0] data_i_3_0[5];
reg valid_i_3_0[5], ready_i_3_0[5];    
wire [`DW-1:0] data_o_3_0[5];
wire valid_o_3_0[5], ready_o_3_0[5];        

reg [`DW-1:0] data_i_3_1[5];
reg valid_i_3_1[5], ready_i_3_1[5];    
wire [`DW-1:0] data_o_3_1[5];
wire valid_o_3_1[5], ready_o_3_1[5];        

reg [`DW-1:0] data_i_3_2[5];
reg valid_i_3_2[5], ready_i_3_2[5];    
wire [`DW-1:0] data_o_3_2[5];
wire valid_o_3_2[5], ready_o_3_2[5];        

reg [`DW-1:0] data_i_3_3[5];
reg valid_i_3_3[5], ready_i_3_3[5];    
wire [`DW-1:0] data_o_3_3[5];
wire valid_o_3_3[5], ready_o_3_3[5];        

reg [`DW-1:0] data_i_3_4[5];
reg valid_i_3_4[5], ready_i_3_4[5];    
wire [`DW-1:0] data_o_3_4[5];
wire valid_o_3_4[5], ready_o_3_4[5];        

reg [`DW-1:0] data_i_3_5[5];
reg valid_i_3_5[5], ready_i_3_5[5];    
wire [`DW-1:0] data_o_3_5[5];
wire valid_o_3_5[5], ready_o_3_5[5];        

reg [`DW-1:0] data_i_3_6[5];
reg valid_i_3_6[5], ready_i_3_6[5];    
wire [`DW-1:0] data_o_3_6[5];
wire valid_o_3_6[5], ready_o_3_6[5];        

reg [`DW-1:0] data_i_3_7[5];
reg valid_i_3_7[5], ready_i_3_7[5];    
wire [`DW-1:0] data_o_3_7[5];
wire valid_o_3_7[5], ready_o_3_7[5];        

reg [`DW-1:0] data_i_3_8[5];
reg valid_i_3_8[5], ready_i_3_8[5];    
wire [`DW-1:0] data_o_3_8[5];
wire valid_o_3_8[5], ready_o_3_8[5];        

reg [`DW-1:0] data_i_3_9[5];
reg valid_i_3_9[5], ready_i_3_9[5];    
wire [`DW-1:0] data_o_3_9[5];
wire valid_o_3_9[5], ready_o_3_9[5];        

reg [`DW-1:0] data_i_3_10[5];
reg valid_i_3_10[5], ready_i_3_10[5];    
wire [`DW-1:0] data_o_3_10[5];
wire valid_o_3_10[5], ready_o_3_10[5];        

reg [`DW-1:0] data_i_3_11[5];
reg valid_i_3_11[5], ready_i_3_11[5];    
wire [`DW-1:0] data_o_3_11[5];
wire valid_o_3_11[5], ready_o_3_11[5];        

reg [`DW-1:0] data_i_3_12[5];
reg valid_i_3_12[5], ready_i_3_12[5];    
wire [`DW-1:0] data_o_3_12[5];
wire valid_o_3_12[5], ready_o_3_12[5];        

reg [`DW-1:0] data_i_3_13[5];
reg valid_i_3_13[5], ready_i_3_13[5];    
wire [`DW-1:0] data_o_3_13[5];
wire valid_o_3_13[5], ready_o_3_13[5];        

reg [`DW-1:0] data_i_3_14[5];
reg valid_i_3_14[5], ready_i_3_14[5];    
wire [`DW-1:0] data_o_3_14[5];
wire valid_o_3_14[5], ready_o_3_14[5];        

reg [`DW-1:0] data_i_3_15[5];
reg valid_i_3_15[5], ready_i_3_15[5];    
wire [`DW-1:0] data_o_3_15[5];
wire valid_o_3_15[5], ready_o_3_15[5];        

reg [`DW-1:0] data_i_3_16[5];
reg valid_i_3_16[5], ready_i_3_16[5];    
wire [`DW-1:0] data_o_3_16[5];
wire valid_o_3_16[5], ready_o_3_16[5];        

reg [`DW-1:0] data_i_3_17[5];
reg valid_i_3_17[5], ready_i_3_17[5];    
wire [`DW-1:0] data_o_3_17[5];
wire valid_o_3_17[5], ready_o_3_17[5];        

reg [`DW-1:0] data_i_3_18[5];
reg valid_i_3_18[5], ready_i_3_18[5];    
wire [`DW-1:0] data_o_3_18[5];
wire valid_o_3_18[5], ready_o_3_18[5];        

reg [`DW-1:0] data_i_3_19[5];
reg valid_i_3_19[5], ready_i_3_19[5];    
wire [`DW-1:0] data_o_3_19[5];
wire valid_o_3_19[5], ready_o_3_19[5];        

reg [`DW-1:0] data_i_3_20[5];
reg valid_i_3_20[5], ready_i_3_20[5];    
wire [`DW-1:0] data_o_3_20[5];
wire valid_o_3_20[5], ready_o_3_20[5];        

reg [`DW-1:0] data_i_3_21[5];
reg valid_i_3_21[5], ready_i_3_21[5];    
wire [`DW-1:0] data_o_3_21[5];
wire valid_o_3_21[5], ready_o_3_21[5];        

reg [`DW-1:0] data_i_3_22[5];
reg valid_i_3_22[5], ready_i_3_22[5];    
wire [`DW-1:0] data_o_3_22[5];
wire valid_o_3_22[5], ready_o_3_22[5];        

reg [`DW-1:0] data_i_3_23[5];
reg valid_i_3_23[5], ready_i_3_23[5];    
wire [`DW-1:0] data_o_3_23[5];
wire valid_o_3_23[5], ready_o_3_23[5];        

reg [`DW-1:0] data_i_3_24[5];
reg valid_i_3_24[5], ready_i_3_24[5];    
wire [`DW-1:0] data_o_3_24[5];
wire valid_o_3_24[5], ready_o_3_24[5];        

reg [`DW-1:0] data_i_4_0[5];
reg valid_i_4_0[5], ready_i_4_0[5];    
wire [`DW-1:0] data_o_4_0[5];
wire valid_o_4_0[5], ready_o_4_0[5];        

reg [`DW-1:0] data_i_4_1[5];
reg valid_i_4_1[5], ready_i_4_1[5];    
wire [`DW-1:0] data_o_4_1[5];
wire valid_o_4_1[5], ready_o_4_1[5];        

reg [`DW-1:0] data_i_4_2[5];
reg valid_i_4_2[5], ready_i_4_2[5];    
wire [`DW-1:0] data_o_4_2[5];
wire valid_o_4_2[5], ready_o_4_2[5];        

reg [`DW-1:0] data_i_4_3[5];
reg valid_i_4_3[5], ready_i_4_3[5];    
wire [`DW-1:0] data_o_4_3[5];
wire valid_o_4_3[5], ready_o_4_3[5];        

reg [`DW-1:0] data_i_4_4[5];
reg valid_i_4_4[5], ready_i_4_4[5];    
wire [`DW-1:0] data_o_4_4[5];
wire valid_o_4_4[5], ready_o_4_4[5];        

reg [`DW-1:0] data_i_4_5[5];
reg valid_i_4_5[5], ready_i_4_5[5];    
wire [`DW-1:0] data_o_4_5[5];
wire valid_o_4_5[5], ready_o_4_5[5];        

reg [`DW-1:0] data_i_4_6[5];
reg valid_i_4_6[5], ready_i_4_6[5];    
wire [`DW-1:0] data_o_4_6[5];
wire valid_o_4_6[5], ready_o_4_6[5];        

reg [`DW-1:0] data_i_4_7[5];
reg valid_i_4_7[5], ready_i_4_7[5];    
wire [`DW-1:0] data_o_4_7[5];
wire valid_o_4_7[5], ready_o_4_7[5];        

reg [`DW-1:0] data_i_4_8[5];
reg valid_i_4_8[5], ready_i_4_8[5];    
wire [`DW-1:0] data_o_4_8[5];
wire valid_o_4_8[5], ready_o_4_8[5];        

reg [`DW-1:0] data_i_4_9[5];
reg valid_i_4_9[5], ready_i_4_9[5];    
wire [`DW-1:0] data_o_4_9[5];
wire valid_o_4_9[5], ready_o_4_9[5];        

reg [`DW-1:0] data_i_4_10[5];
reg valid_i_4_10[5], ready_i_4_10[5];    
wire [`DW-1:0] data_o_4_10[5];
wire valid_o_4_10[5], ready_o_4_10[5];        

reg [`DW-1:0] data_i_4_11[5];
reg valid_i_4_11[5], ready_i_4_11[5];    
wire [`DW-1:0] data_o_4_11[5];
wire valid_o_4_11[5], ready_o_4_11[5];        

reg [`DW-1:0] data_i_4_12[5];
reg valid_i_4_12[5], ready_i_4_12[5];    
wire [`DW-1:0] data_o_4_12[5];
wire valid_o_4_12[5], ready_o_4_12[5];        

reg [`DW-1:0] data_i_4_13[5];
reg valid_i_4_13[5], ready_i_4_13[5];    
wire [`DW-1:0] data_o_4_13[5];
wire valid_o_4_13[5], ready_o_4_13[5];        

reg [`DW-1:0] data_i_4_14[5];
reg valid_i_4_14[5], ready_i_4_14[5];    
wire [`DW-1:0] data_o_4_14[5];
wire valid_o_4_14[5], ready_o_4_14[5];        

reg [`DW-1:0] data_i_4_15[5];
reg valid_i_4_15[5], ready_i_4_15[5];    
wire [`DW-1:0] data_o_4_15[5];
wire valid_o_4_15[5], ready_o_4_15[5];        

reg [`DW-1:0] data_i_4_16[5];
reg valid_i_4_16[5], ready_i_4_16[5];    
wire [`DW-1:0] data_o_4_16[5];
wire valid_o_4_16[5], ready_o_4_16[5];        

reg [`DW-1:0] data_i_4_17[5];
reg valid_i_4_17[5], ready_i_4_17[5];    
wire [`DW-1:0] data_o_4_17[5];
wire valid_o_4_17[5], ready_o_4_17[5];        

reg [`DW-1:0] data_i_4_18[5];
reg valid_i_4_18[5], ready_i_4_18[5];    
wire [`DW-1:0] data_o_4_18[5];
wire valid_o_4_18[5], ready_o_4_18[5];        

reg [`DW-1:0] data_i_4_19[5];
reg valid_i_4_19[5], ready_i_4_19[5];    
wire [`DW-1:0] data_o_4_19[5];
wire valid_o_4_19[5], ready_o_4_19[5];        

reg [`DW-1:0] data_i_4_20[5];
reg valid_i_4_20[5], ready_i_4_20[5];    
wire [`DW-1:0] data_o_4_20[5];
wire valid_o_4_20[5], ready_o_4_20[5];        

reg [`DW-1:0] data_i_4_21[5];
reg valid_i_4_21[5], ready_i_4_21[5];    
wire [`DW-1:0] data_o_4_21[5];
wire valid_o_4_21[5], ready_o_4_21[5];        

reg [`DW-1:0] data_i_4_22[5];
reg valid_i_4_22[5], ready_i_4_22[5];    
wire [`DW-1:0] data_o_4_22[5];
wire valid_o_4_22[5], ready_o_4_22[5];        

reg [`DW-1:0] data_i_4_23[5];
reg valid_i_4_23[5], ready_i_4_23[5];    
wire [`DW-1:0] data_o_4_23[5];
wire valid_o_4_23[5], ready_o_4_23[5];        

reg [`DW-1:0] data_i_4_24[5];
reg valid_i_4_24[5], ready_i_4_24[5];    
wire [`DW-1:0] data_o_4_24[5];
wire valid_o_4_24[5], ready_o_4_24[5];        

reg [`DW-1:0] data_i_5_0[5];
reg valid_i_5_0[5], ready_i_5_0[5];    
wire [`DW-1:0] data_o_5_0[5];
wire valid_o_5_0[5], ready_o_5_0[5];        

reg [`DW-1:0] data_i_5_1[5];
reg valid_i_5_1[5], ready_i_5_1[5];    
wire [`DW-1:0] data_o_5_1[5];
wire valid_o_5_1[5], ready_o_5_1[5];        

reg [`DW-1:0] data_i_5_2[5];
reg valid_i_5_2[5], ready_i_5_2[5];    
wire [`DW-1:0] data_o_5_2[5];
wire valid_o_5_2[5], ready_o_5_2[5];        

reg [`DW-1:0] data_i_5_3[5];
reg valid_i_5_3[5], ready_i_5_3[5];    
wire [`DW-1:0] data_o_5_3[5];
wire valid_o_5_3[5], ready_o_5_3[5];        

reg [`DW-1:0] data_i_5_4[5];
reg valid_i_5_4[5], ready_i_5_4[5];    
wire [`DW-1:0] data_o_5_4[5];
wire valid_o_5_4[5], ready_o_5_4[5];        

reg [`DW-1:0] data_i_5_5[5];
reg valid_i_5_5[5], ready_i_5_5[5];    
wire [`DW-1:0] data_o_5_5[5];
wire valid_o_5_5[5], ready_o_5_5[5];        

reg [`DW-1:0] data_i_5_6[5];
reg valid_i_5_6[5], ready_i_5_6[5];    
wire [`DW-1:0] data_o_5_6[5];
wire valid_o_5_6[5], ready_o_5_6[5];        

reg [`DW-1:0] data_i_5_7[5];
reg valid_i_5_7[5], ready_i_5_7[5];    
wire [`DW-1:0] data_o_5_7[5];
wire valid_o_5_7[5], ready_o_5_7[5];        

reg [`DW-1:0] data_i_5_8[5];
reg valid_i_5_8[5], ready_i_5_8[5];    
wire [`DW-1:0] data_o_5_8[5];
wire valid_o_5_8[5], ready_o_5_8[5];        

reg [`DW-1:0] data_i_5_9[5];
reg valid_i_5_9[5], ready_i_5_9[5];    
wire [`DW-1:0] data_o_5_9[5];
wire valid_o_5_9[5], ready_o_5_9[5];        

reg [`DW-1:0] data_i_5_10[5];
reg valid_i_5_10[5], ready_i_5_10[5];    
wire [`DW-1:0] data_o_5_10[5];
wire valid_o_5_10[5], ready_o_5_10[5];        

reg [`DW-1:0] data_i_5_11[5];
reg valid_i_5_11[5], ready_i_5_11[5];    
wire [`DW-1:0] data_o_5_11[5];
wire valid_o_5_11[5], ready_o_5_11[5];        

reg [`DW-1:0] data_i_5_12[5];
reg valid_i_5_12[5], ready_i_5_12[5];    
wire [`DW-1:0] data_o_5_12[5];
wire valid_o_5_12[5], ready_o_5_12[5];        

reg [`DW-1:0] data_i_5_13[5];
reg valid_i_5_13[5], ready_i_5_13[5];    
wire [`DW-1:0] data_o_5_13[5];
wire valid_o_5_13[5], ready_o_5_13[5];        

reg [`DW-1:0] data_i_5_14[5];
reg valid_i_5_14[5], ready_i_5_14[5];    
wire [`DW-1:0] data_o_5_14[5];
wire valid_o_5_14[5], ready_o_5_14[5];        

reg [`DW-1:0] data_i_5_15[5];
reg valid_i_5_15[5], ready_i_5_15[5];    
wire [`DW-1:0] data_o_5_15[5];
wire valid_o_5_15[5], ready_o_5_15[5];        

reg [`DW-1:0] data_i_5_16[5];
reg valid_i_5_16[5], ready_i_5_16[5];    
wire [`DW-1:0] data_o_5_16[5];
wire valid_o_5_16[5], ready_o_5_16[5];        

reg [`DW-1:0] data_i_5_17[5];
reg valid_i_5_17[5], ready_i_5_17[5];    
wire [`DW-1:0] data_o_5_17[5];
wire valid_o_5_17[5], ready_o_5_17[5];        

reg [`DW-1:0] data_i_5_18[5];
reg valid_i_5_18[5], ready_i_5_18[5];    
wire [`DW-1:0] data_o_5_18[5];
wire valid_o_5_18[5], ready_o_5_18[5];        

reg [`DW-1:0] data_i_5_19[5];
reg valid_i_5_19[5], ready_i_5_19[5];    
wire [`DW-1:0] data_o_5_19[5];
wire valid_o_5_19[5], ready_o_5_19[5];        

reg [`DW-1:0] data_i_5_20[5];
reg valid_i_5_20[5], ready_i_5_20[5];    
wire [`DW-1:0] data_o_5_20[5];
wire valid_o_5_20[5], ready_o_5_20[5];        

reg [`DW-1:0] data_i_5_21[5];
reg valid_i_5_21[5], ready_i_5_21[5];    
wire [`DW-1:0] data_o_5_21[5];
wire valid_o_5_21[5], ready_o_5_21[5];        

reg [`DW-1:0] data_i_5_22[5];
reg valid_i_5_22[5], ready_i_5_22[5];    
wire [`DW-1:0] data_o_5_22[5];
wire valid_o_5_22[5], ready_o_5_22[5];        

reg [`DW-1:0] data_i_5_23[5];
reg valid_i_5_23[5], ready_i_5_23[5];    
wire [`DW-1:0] data_o_5_23[5];
wire valid_o_5_23[5], ready_o_5_23[5];        

reg [`DW-1:0] data_i_5_24[5];
reg valid_i_5_24[5], ready_i_5_24[5];    
wire [`DW-1:0] data_o_5_24[5];
wire valid_o_5_24[5], ready_o_5_24[5];        

reg [`DW-1:0] data_i_6_0[5];
reg valid_i_6_0[5], ready_i_6_0[5];    
wire [`DW-1:0] data_o_6_0[5];
wire valid_o_6_0[5], ready_o_6_0[5];        

reg [`DW-1:0] data_i_6_1[5];
reg valid_i_6_1[5], ready_i_6_1[5];    
wire [`DW-1:0] data_o_6_1[5];
wire valid_o_6_1[5], ready_o_6_1[5];        

reg [`DW-1:0] data_i_6_2[5];
reg valid_i_6_2[5], ready_i_6_2[5];    
wire [`DW-1:0] data_o_6_2[5];
wire valid_o_6_2[5], ready_o_6_2[5];        

reg [`DW-1:0] data_i_6_3[5];
reg valid_i_6_3[5], ready_i_6_3[5];    
wire [`DW-1:0] data_o_6_3[5];
wire valid_o_6_3[5], ready_o_6_3[5];        

reg [`DW-1:0] data_i_6_4[5];
reg valid_i_6_4[5], ready_i_6_4[5];    
wire [`DW-1:0] data_o_6_4[5];
wire valid_o_6_4[5], ready_o_6_4[5];        

reg [`DW-1:0] data_i_6_5[5];
reg valid_i_6_5[5], ready_i_6_5[5];    
wire [`DW-1:0] data_o_6_5[5];
wire valid_o_6_5[5], ready_o_6_5[5];        

reg [`DW-1:0] data_i_6_6[5];
reg valid_i_6_6[5], ready_i_6_6[5];    
wire [`DW-1:0] data_o_6_6[5];
wire valid_o_6_6[5], ready_o_6_6[5];        

reg [`DW-1:0] data_i_6_7[5];
reg valid_i_6_7[5], ready_i_6_7[5];    
wire [`DW-1:0] data_o_6_7[5];
wire valid_o_6_7[5], ready_o_6_7[5];        

reg [`DW-1:0] data_i_6_8[5];
reg valid_i_6_8[5], ready_i_6_8[5];    
wire [`DW-1:0] data_o_6_8[5];
wire valid_o_6_8[5], ready_o_6_8[5];        

reg [`DW-1:0] data_i_6_9[5];
reg valid_i_6_9[5], ready_i_6_9[5];    
wire [`DW-1:0] data_o_6_9[5];
wire valid_o_6_9[5], ready_o_6_9[5];        

reg [`DW-1:0] data_i_6_10[5];
reg valid_i_6_10[5], ready_i_6_10[5];    
wire [`DW-1:0] data_o_6_10[5];
wire valid_o_6_10[5], ready_o_6_10[5];        

reg [`DW-1:0] data_i_6_11[5];
reg valid_i_6_11[5], ready_i_6_11[5];    
wire [`DW-1:0] data_o_6_11[5];
wire valid_o_6_11[5], ready_o_6_11[5];        

reg [`DW-1:0] data_i_6_12[5];
reg valid_i_6_12[5], ready_i_6_12[5];    
wire [`DW-1:0] data_o_6_12[5];
wire valid_o_6_12[5], ready_o_6_12[5];        

reg [`DW-1:0] data_i_6_13[5];
reg valid_i_6_13[5], ready_i_6_13[5];    
wire [`DW-1:0] data_o_6_13[5];
wire valid_o_6_13[5], ready_o_6_13[5];        

reg [`DW-1:0] data_i_6_14[5];
reg valid_i_6_14[5], ready_i_6_14[5];    
wire [`DW-1:0] data_o_6_14[5];
wire valid_o_6_14[5], ready_o_6_14[5];        

reg [`DW-1:0] data_i_6_15[5];
reg valid_i_6_15[5], ready_i_6_15[5];    
wire [`DW-1:0] data_o_6_15[5];
wire valid_o_6_15[5], ready_o_6_15[5];        

reg [`DW-1:0] data_i_6_16[5];
reg valid_i_6_16[5], ready_i_6_16[5];    
wire [`DW-1:0] data_o_6_16[5];
wire valid_o_6_16[5], ready_o_6_16[5];        

reg [`DW-1:0] data_i_6_17[5];
reg valid_i_6_17[5], ready_i_6_17[5];    
wire [`DW-1:0] data_o_6_17[5];
wire valid_o_6_17[5], ready_o_6_17[5];        

reg [`DW-1:0] data_i_6_18[5];
reg valid_i_6_18[5], ready_i_6_18[5];    
wire [`DW-1:0] data_o_6_18[5];
wire valid_o_6_18[5], ready_o_6_18[5];        

reg [`DW-1:0] data_i_6_19[5];
reg valid_i_6_19[5], ready_i_6_19[5];    
wire [`DW-1:0] data_o_6_19[5];
wire valid_o_6_19[5], ready_o_6_19[5];        

reg [`DW-1:0] data_i_6_20[5];
reg valid_i_6_20[5], ready_i_6_20[5];    
wire [`DW-1:0] data_o_6_20[5];
wire valid_o_6_20[5], ready_o_6_20[5];        

reg [`DW-1:0] data_i_6_21[5];
reg valid_i_6_21[5], ready_i_6_21[5];    
wire [`DW-1:0] data_o_6_21[5];
wire valid_o_6_21[5], ready_o_6_21[5];        

reg [`DW-1:0] data_i_6_22[5];
reg valid_i_6_22[5], ready_i_6_22[5];    
wire [`DW-1:0] data_o_6_22[5];
wire valid_o_6_22[5], ready_o_6_22[5];        

reg [`DW-1:0] data_i_6_23[5];
reg valid_i_6_23[5], ready_i_6_23[5];    
wire [`DW-1:0] data_o_6_23[5];
wire valid_o_6_23[5], ready_o_6_23[5];        

reg [`DW-1:0] data_i_6_24[5];
reg valid_i_6_24[5], ready_i_6_24[5];    
wire [`DW-1:0] data_o_6_24[5];
wire valid_o_6_24[5], ready_o_6_24[5];        

reg [`DW-1:0] data_i_7_0[5];
reg valid_i_7_0[5], ready_i_7_0[5];    
wire [`DW-1:0] data_o_7_0[5];
wire valid_o_7_0[5], ready_o_7_0[5];        

reg [`DW-1:0] data_i_7_1[5];
reg valid_i_7_1[5], ready_i_7_1[5];    
wire [`DW-1:0] data_o_7_1[5];
wire valid_o_7_1[5], ready_o_7_1[5];        

reg [`DW-1:0] data_i_7_2[5];
reg valid_i_7_2[5], ready_i_7_2[5];    
wire [`DW-1:0] data_o_7_2[5];
wire valid_o_7_2[5], ready_o_7_2[5];        

reg [`DW-1:0] data_i_7_3[5];
reg valid_i_7_3[5], ready_i_7_3[5];    
wire [`DW-1:0] data_o_7_3[5];
wire valid_o_7_3[5], ready_o_7_3[5];        

reg [`DW-1:0] data_i_7_4[5];
reg valid_i_7_4[5], ready_i_7_4[5];    
wire [`DW-1:0] data_o_7_4[5];
wire valid_o_7_4[5], ready_o_7_4[5];        

reg [`DW-1:0] data_i_7_5[5];
reg valid_i_7_5[5], ready_i_7_5[5];    
wire [`DW-1:0] data_o_7_5[5];
wire valid_o_7_5[5], ready_o_7_5[5];        

reg [`DW-1:0] data_i_7_6[5];
reg valid_i_7_6[5], ready_i_7_6[5];    
wire [`DW-1:0] data_o_7_6[5];
wire valid_o_7_6[5], ready_o_7_6[5];        

reg [`DW-1:0] data_i_7_7[5];
reg valid_i_7_7[5], ready_i_7_7[5];    
wire [`DW-1:0] data_o_7_7[5];
wire valid_o_7_7[5], ready_o_7_7[5];        

reg [`DW-1:0] data_i_7_8[5];
reg valid_i_7_8[5], ready_i_7_8[5];    
wire [`DW-1:0] data_o_7_8[5];
wire valid_o_7_8[5], ready_o_7_8[5];        

reg [`DW-1:0] data_i_7_9[5];
reg valid_i_7_9[5], ready_i_7_9[5];    
wire [`DW-1:0] data_o_7_9[5];
wire valid_o_7_9[5], ready_o_7_9[5];        

reg [`DW-1:0] data_i_7_10[5];
reg valid_i_7_10[5], ready_i_7_10[5];    
wire [`DW-1:0] data_o_7_10[5];
wire valid_o_7_10[5], ready_o_7_10[5];        

reg [`DW-1:0] data_i_7_11[5];
reg valid_i_7_11[5], ready_i_7_11[5];    
wire [`DW-1:0] data_o_7_11[5];
wire valid_o_7_11[5], ready_o_7_11[5];        

reg [`DW-1:0] data_i_7_12[5];
reg valid_i_7_12[5], ready_i_7_12[5];    
wire [`DW-1:0] data_o_7_12[5];
wire valid_o_7_12[5], ready_o_7_12[5];        

reg [`DW-1:0] data_i_7_13[5];
reg valid_i_7_13[5], ready_i_7_13[5];    
wire [`DW-1:0] data_o_7_13[5];
wire valid_o_7_13[5], ready_o_7_13[5];        

reg [`DW-1:0] data_i_7_14[5];
reg valid_i_7_14[5], ready_i_7_14[5];    
wire [`DW-1:0] data_o_7_14[5];
wire valid_o_7_14[5], ready_o_7_14[5];        

reg [`DW-1:0] data_i_7_15[5];
reg valid_i_7_15[5], ready_i_7_15[5];    
wire [`DW-1:0] data_o_7_15[5];
wire valid_o_7_15[5], ready_o_7_15[5];        

reg [`DW-1:0] data_i_7_16[5];
reg valid_i_7_16[5], ready_i_7_16[5];    
wire [`DW-1:0] data_o_7_16[5];
wire valid_o_7_16[5], ready_o_7_16[5];        

reg [`DW-1:0] data_i_7_17[5];
reg valid_i_7_17[5], ready_i_7_17[5];    
wire [`DW-1:0] data_o_7_17[5];
wire valid_o_7_17[5], ready_o_7_17[5];        

reg [`DW-1:0] data_i_7_18[5];
reg valid_i_7_18[5], ready_i_7_18[5];    
wire [`DW-1:0] data_o_7_18[5];
wire valid_o_7_18[5], ready_o_7_18[5];        

reg [`DW-1:0] data_i_7_19[5];
reg valid_i_7_19[5], ready_i_7_19[5];    
wire [`DW-1:0] data_o_7_19[5];
wire valid_o_7_19[5], ready_o_7_19[5];        

reg [`DW-1:0] data_i_7_20[5];
reg valid_i_7_20[5], ready_i_7_20[5];    
wire [`DW-1:0] data_o_7_20[5];
wire valid_o_7_20[5], ready_o_7_20[5];        

reg [`DW-1:0] data_i_7_21[5];
reg valid_i_7_21[5], ready_i_7_21[5];    
wire [`DW-1:0] data_o_7_21[5];
wire valid_o_7_21[5], ready_o_7_21[5];        

reg [`DW-1:0] data_i_7_22[5];
reg valid_i_7_22[5], ready_i_7_22[5];    
wire [`DW-1:0] data_o_7_22[5];
wire valid_o_7_22[5], ready_o_7_22[5];        

reg [`DW-1:0] data_i_7_23[5];
reg valid_i_7_23[5], ready_i_7_23[5];    
wire [`DW-1:0] data_o_7_23[5];
wire valid_o_7_23[5], ready_o_7_23[5];        

reg [`DW-1:0] data_i_7_24[5];
reg valid_i_7_24[5], ready_i_7_24[5];    
wire [`DW-1:0] data_o_7_24[5];
wire valid_o_7_24[5], ready_o_7_24[5];        

reg [`DW-1:0] data_i_8_0[5];
reg valid_i_8_0[5], ready_i_8_0[5];    
wire [`DW-1:0] data_o_8_0[5];
wire valid_o_8_0[5], ready_o_8_0[5];        

reg [`DW-1:0] data_i_8_1[5];
reg valid_i_8_1[5], ready_i_8_1[5];    
wire [`DW-1:0] data_o_8_1[5];
wire valid_o_8_1[5], ready_o_8_1[5];        

reg [`DW-1:0] data_i_8_2[5];
reg valid_i_8_2[5], ready_i_8_2[5];    
wire [`DW-1:0] data_o_8_2[5];
wire valid_o_8_2[5], ready_o_8_2[5];        

reg [`DW-1:0] data_i_8_3[5];
reg valid_i_8_3[5], ready_i_8_3[5];    
wire [`DW-1:0] data_o_8_3[5];
wire valid_o_8_3[5], ready_o_8_3[5];        

reg [`DW-1:0] data_i_8_4[5];
reg valid_i_8_4[5], ready_i_8_4[5];    
wire [`DW-1:0] data_o_8_4[5];
wire valid_o_8_4[5], ready_o_8_4[5];        

reg [`DW-1:0] data_i_8_5[5];
reg valid_i_8_5[5], ready_i_8_5[5];    
wire [`DW-1:0] data_o_8_5[5];
wire valid_o_8_5[5], ready_o_8_5[5];        

reg [`DW-1:0] data_i_8_6[5];
reg valid_i_8_6[5], ready_i_8_6[5];    
wire [`DW-1:0] data_o_8_6[5];
wire valid_o_8_6[5], ready_o_8_6[5];        

reg [`DW-1:0] data_i_8_7[5];
reg valid_i_8_7[5], ready_i_8_7[5];    
wire [`DW-1:0] data_o_8_7[5];
wire valid_o_8_7[5], ready_o_8_7[5];        

reg [`DW-1:0] data_i_8_8[5];
reg valid_i_8_8[5], ready_i_8_8[5];    
wire [`DW-1:0] data_o_8_8[5];
wire valid_o_8_8[5], ready_o_8_8[5];        

reg [`DW-1:0] data_i_8_9[5];
reg valid_i_8_9[5], ready_i_8_9[5];    
wire [`DW-1:0] data_o_8_9[5];
wire valid_o_8_9[5], ready_o_8_9[5];        

reg [`DW-1:0] data_i_8_10[5];
reg valid_i_8_10[5], ready_i_8_10[5];    
wire [`DW-1:0] data_o_8_10[5];
wire valid_o_8_10[5], ready_o_8_10[5];        

reg [`DW-1:0] data_i_8_11[5];
reg valid_i_8_11[5], ready_i_8_11[5];    
wire [`DW-1:0] data_o_8_11[5];
wire valid_o_8_11[5], ready_o_8_11[5];        

reg [`DW-1:0] data_i_8_12[5];
reg valid_i_8_12[5], ready_i_8_12[5];    
wire [`DW-1:0] data_o_8_12[5];
wire valid_o_8_12[5], ready_o_8_12[5];        

reg [`DW-1:0] data_i_8_13[5];
reg valid_i_8_13[5], ready_i_8_13[5];    
wire [`DW-1:0] data_o_8_13[5];
wire valid_o_8_13[5], ready_o_8_13[5];        

reg [`DW-1:0] data_i_8_14[5];
reg valid_i_8_14[5], ready_i_8_14[5];    
wire [`DW-1:0] data_o_8_14[5];
wire valid_o_8_14[5], ready_o_8_14[5];        

reg [`DW-1:0] data_i_8_15[5];
reg valid_i_8_15[5], ready_i_8_15[5];    
wire [`DW-1:0] data_o_8_15[5];
wire valid_o_8_15[5], ready_o_8_15[5];        

reg [`DW-1:0] data_i_8_16[5];
reg valid_i_8_16[5], ready_i_8_16[5];    
wire [`DW-1:0] data_o_8_16[5];
wire valid_o_8_16[5], ready_o_8_16[5];        

reg [`DW-1:0] data_i_8_17[5];
reg valid_i_8_17[5], ready_i_8_17[5];    
wire [`DW-1:0] data_o_8_17[5];
wire valid_o_8_17[5], ready_o_8_17[5];        

reg [`DW-1:0] data_i_8_18[5];
reg valid_i_8_18[5], ready_i_8_18[5];    
wire [`DW-1:0] data_o_8_18[5];
wire valid_o_8_18[5], ready_o_8_18[5];        

reg [`DW-1:0] data_i_8_19[5];
reg valid_i_8_19[5], ready_i_8_19[5];    
wire [`DW-1:0] data_o_8_19[5];
wire valid_o_8_19[5], ready_o_8_19[5];        

reg [`DW-1:0] data_i_8_20[5];
reg valid_i_8_20[5], ready_i_8_20[5];    
wire [`DW-1:0] data_o_8_20[5];
wire valid_o_8_20[5], ready_o_8_20[5];        

reg [`DW-1:0] data_i_8_21[5];
reg valid_i_8_21[5], ready_i_8_21[5];    
wire [`DW-1:0] data_o_8_21[5];
wire valid_o_8_21[5], ready_o_8_21[5];        

reg [`DW-1:0] data_i_8_22[5];
reg valid_i_8_22[5], ready_i_8_22[5];    
wire [`DW-1:0] data_o_8_22[5];
wire valid_o_8_22[5], ready_o_8_22[5];        

reg [`DW-1:0] data_i_8_23[5];
reg valid_i_8_23[5], ready_i_8_23[5];    
wire [`DW-1:0] data_o_8_23[5];
wire valid_o_8_23[5], ready_o_8_23[5];        

reg [`DW-1:0] data_i_8_24[5];
reg valid_i_8_24[5], ready_i_8_24[5];    
wire [`DW-1:0] data_o_8_24[5];
wire valid_o_8_24[5], ready_o_8_24[5];        

reg [`DW-1:0] data_i_9_0[5];
reg valid_i_9_0[5], ready_i_9_0[5];    
wire [`DW-1:0] data_o_9_0[5];
wire valid_o_9_0[5], ready_o_9_0[5];        

reg [`DW-1:0] data_i_9_1[5];
reg valid_i_9_1[5], ready_i_9_1[5];    
wire [`DW-1:0] data_o_9_1[5];
wire valid_o_9_1[5], ready_o_9_1[5];        

reg [`DW-1:0] data_i_9_2[5];
reg valid_i_9_2[5], ready_i_9_2[5];    
wire [`DW-1:0] data_o_9_2[5];
wire valid_o_9_2[5], ready_o_9_2[5];        

reg [`DW-1:0] data_i_9_3[5];
reg valid_i_9_3[5], ready_i_9_3[5];    
wire [`DW-1:0] data_o_9_3[5];
wire valid_o_9_3[5], ready_o_9_3[5];        

reg [`DW-1:0] data_i_9_4[5];
reg valid_i_9_4[5], ready_i_9_4[5];    
wire [`DW-1:0] data_o_9_4[5];
wire valid_o_9_4[5], ready_o_9_4[5];        

reg [`DW-1:0] data_i_9_5[5];
reg valid_i_9_5[5], ready_i_9_5[5];    
wire [`DW-1:0] data_o_9_5[5];
wire valid_o_9_5[5], ready_o_9_5[5];        

reg [`DW-1:0] data_i_9_6[5];
reg valid_i_9_6[5], ready_i_9_6[5];    
wire [`DW-1:0] data_o_9_6[5];
wire valid_o_9_6[5], ready_o_9_6[5];        

reg [`DW-1:0] data_i_9_7[5];
reg valid_i_9_7[5], ready_i_9_7[5];    
wire [`DW-1:0] data_o_9_7[5];
wire valid_o_9_7[5], ready_o_9_7[5];        

reg [`DW-1:0] data_i_9_8[5];
reg valid_i_9_8[5], ready_i_9_8[5];    
wire [`DW-1:0] data_o_9_8[5];
wire valid_o_9_8[5], ready_o_9_8[5];        

reg [`DW-1:0] data_i_9_9[5];
reg valid_i_9_9[5], ready_i_9_9[5];    
wire [`DW-1:0] data_o_9_9[5];
wire valid_o_9_9[5], ready_o_9_9[5];        

reg [`DW-1:0] data_i_9_10[5];
reg valid_i_9_10[5], ready_i_9_10[5];    
wire [`DW-1:0] data_o_9_10[5];
wire valid_o_9_10[5], ready_o_9_10[5];        

reg [`DW-1:0] data_i_9_11[5];
reg valid_i_9_11[5], ready_i_9_11[5];    
wire [`DW-1:0] data_o_9_11[5];
wire valid_o_9_11[5], ready_o_9_11[5];        

reg [`DW-1:0] data_i_9_12[5];
reg valid_i_9_12[5], ready_i_9_12[5];    
wire [`DW-1:0] data_o_9_12[5];
wire valid_o_9_12[5], ready_o_9_12[5];        

reg [`DW-1:0] data_i_9_13[5];
reg valid_i_9_13[5], ready_i_9_13[5];    
wire [`DW-1:0] data_o_9_13[5];
wire valid_o_9_13[5], ready_o_9_13[5];        

reg [`DW-1:0] data_i_9_14[5];
reg valid_i_9_14[5], ready_i_9_14[5];    
wire [`DW-1:0] data_o_9_14[5];
wire valid_o_9_14[5], ready_o_9_14[5];        

reg [`DW-1:0] data_i_9_15[5];
reg valid_i_9_15[5], ready_i_9_15[5];    
wire [`DW-1:0] data_o_9_15[5];
wire valid_o_9_15[5], ready_o_9_15[5];        

reg [`DW-1:0] data_i_9_16[5];
reg valid_i_9_16[5], ready_i_9_16[5];    
wire [`DW-1:0] data_o_9_16[5];
wire valid_o_9_16[5], ready_o_9_16[5];        

reg [`DW-1:0] data_i_9_17[5];
reg valid_i_9_17[5], ready_i_9_17[5];    
wire [`DW-1:0] data_o_9_17[5];
wire valid_o_9_17[5], ready_o_9_17[5];        

reg [`DW-1:0] data_i_9_18[5];
reg valid_i_9_18[5], ready_i_9_18[5];    
wire [`DW-1:0] data_o_9_18[5];
wire valid_o_9_18[5], ready_o_9_18[5];        

reg [`DW-1:0] data_i_9_19[5];
reg valid_i_9_19[5], ready_i_9_19[5];    
wire [`DW-1:0] data_o_9_19[5];
wire valid_o_9_19[5], ready_o_9_19[5];        

reg [`DW-1:0] data_i_9_20[5];
reg valid_i_9_20[5], ready_i_9_20[5];    
wire [`DW-1:0] data_o_9_20[5];
wire valid_o_9_20[5], ready_o_9_20[5];        

reg [`DW-1:0] data_i_9_21[5];
reg valid_i_9_21[5], ready_i_9_21[5];    
wire [`DW-1:0] data_o_9_21[5];
wire valid_o_9_21[5], ready_o_9_21[5];        

reg [`DW-1:0] data_i_9_22[5];
reg valid_i_9_22[5], ready_i_9_22[5];    
wire [`DW-1:0] data_o_9_22[5];
wire valid_o_9_22[5], ready_o_9_22[5];        

reg [`DW-1:0] data_i_9_23[5];
reg valid_i_9_23[5], ready_i_9_23[5];    
wire [`DW-1:0] data_o_9_23[5];
wire valid_o_9_23[5], ready_o_9_23[5];        

reg [`DW-1:0] data_i_9_24[5];
reg valid_i_9_24[5], ready_i_9_24[5];    
wire [`DW-1:0] data_o_9_24[5];
wire valid_o_9_24[5], ready_o_9_24[5];        

always@(*) begin
    data_o[0][0] = data_o_0_0[0];
    valid_o[0][0] = valid_o_0_0[0];
    ready_o[0][0] = ready_o_0_0[0];
    data_o[0][1] = data_o_0_1[0];
    valid_o[0][1] = valid_o_0_1[0];
    ready_o[0][1] = ready_o_0_1[0];
    data_o[0][2] = data_o_0_2[0];
    valid_o[0][2] = valid_o_0_2[0];
    ready_o[0][2] = ready_o_0_2[0];
    data_o[0][3] = data_o_0_3[0];
    valid_o[0][3] = valid_o_0_3[0];
    ready_o[0][3] = ready_o_0_3[0];
    data_o[0][4] = data_o_0_4[0];
    valid_o[0][4] = valid_o_0_4[0];
    ready_o[0][4] = ready_o_0_4[0];
    data_o[0][5] = data_o_0_5[0];
    valid_o[0][5] = valid_o_0_5[0];
    ready_o[0][5] = ready_o_0_5[0];
    data_o[0][6] = data_o_0_6[0];
    valid_o[0][6] = valid_o_0_6[0];
    ready_o[0][6] = ready_o_0_6[0];
    data_o[0][7] = data_o_0_7[0];
    valid_o[0][7] = valid_o_0_7[0];
    ready_o[0][7] = ready_o_0_7[0];
    data_o[0][8] = data_o_0_8[0];
    valid_o[0][8] = valid_o_0_8[0];
    ready_o[0][8] = ready_o_0_8[0];
    data_o[0][9] = data_o_0_9[0];
    valid_o[0][9] = valid_o_0_9[0];
    ready_o[0][9] = ready_o_0_9[0];
    data_o[0][10] = data_o_0_10[0];
    valid_o[0][10] = valid_o_0_10[0];
    ready_o[0][10] = ready_o_0_10[0];
    data_o[0][11] = data_o_0_11[0];
    valid_o[0][11] = valid_o_0_11[0];
    ready_o[0][11] = ready_o_0_11[0];
    data_o[0][12] = data_o_0_12[0];
    valid_o[0][12] = valid_o_0_12[0];
    ready_o[0][12] = ready_o_0_12[0];
    data_o[0][13] = data_o_0_13[0];
    valid_o[0][13] = valid_o_0_13[0];
    ready_o[0][13] = ready_o_0_13[0];
    data_o[0][14] = data_o_0_14[0];
    valid_o[0][14] = valid_o_0_14[0];
    ready_o[0][14] = ready_o_0_14[0];
    data_o[0][15] = data_o_0_15[0];
    valid_o[0][15] = valid_o_0_15[0];
    ready_o[0][15] = ready_o_0_15[0];
    data_o[0][16] = data_o_0_16[0];
    valid_o[0][16] = valid_o_0_16[0];
    ready_o[0][16] = ready_o_0_16[0];
    data_o[0][17] = data_o_0_17[0];
    valid_o[0][17] = valid_o_0_17[0];
    ready_o[0][17] = ready_o_0_17[0];
    data_o[0][18] = data_o_0_18[0];
    valid_o[0][18] = valid_o_0_18[0];
    ready_o[0][18] = ready_o_0_18[0];
    data_o[0][19] = data_o_0_19[0];
    valid_o[0][19] = valid_o_0_19[0];
    ready_o[0][19] = ready_o_0_19[0];
    data_o[0][20] = data_o_0_20[0];
    valid_o[0][20] = valid_o_0_20[0];
    ready_o[0][20] = ready_o_0_20[0];
    data_o[0][21] = data_o_0_21[0];
    valid_o[0][21] = valid_o_0_21[0];
    ready_o[0][21] = ready_o_0_21[0];
    data_o[0][22] = data_o_0_22[0];
    valid_o[0][22] = valid_o_0_22[0];
    ready_o[0][22] = ready_o_0_22[0];
    data_o[0][23] = data_o_0_23[0];
    valid_o[0][23] = valid_o_0_23[0];
    ready_o[0][23] = ready_o_0_23[0];
    data_o[0][24] = data_o_0_24[0];
    valid_o[0][24] = valid_o_0_24[0];
    ready_o[0][24] = ready_o_0_24[0];
    data_o[1][0] = data_o_1_0[0];
    valid_o[1][0] = valid_o_1_0[0];
    ready_o[1][0] = ready_o_1_0[0];
    data_o[1][1] = data_o_1_1[0];
    valid_o[1][1] = valid_o_1_1[0];
    ready_o[1][1] = ready_o_1_1[0];
    data_o[1][2] = data_o_1_2[0];
    valid_o[1][2] = valid_o_1_2[0];
    ready_o[1][2] = ready_o_1_2[0];
    data_o[1][3] = data_o_1_3[0];
    valid_o[1][3] = valid_o_1_3[0];
    ready_o[1][3] = ready_o_1_3[0];
    data_o[1][4] = data_o_1_4[0];
    valid_o[1][4] = valid_o_1_4[0];
    ready_o[1][4] = ready_o_1_4[0];
    data_o[1][5] = data_o_1_5[0];
    valid_o[1][5] = valid_o_1_5[0];
    ready_o[1][5] = ready_o_1_5[0];
    data_o[1][6] = data_o_1_6[0];
    valid_o[1][6] = valid_o_1_6[0];
    ready_o[1][6] = ready_o_1_6[0];
    data_o[1][7] = data_o_1_7[0];
    valid_o[1][7] = valid_o_1_7[0];
    ready_o[1][7] = ready_o_1_7[0];
    data_o[1][8] = data_o_1_8[0];
    valid_o[1][8] = valid_o_1_8[0];
    ready_o[1][8] = ready_o_1_8[0];
    data_o[1][9] = data_o_1_9[0];
    valid_o[1][9] = valid_o_1_9[0];
    ready_o[1][9] = ready_o_1_9[0];
    data_o[1][10] = data_o_1_10[0];
    valid_o[1][10] = valid_o_1_10[0];
    ready_o[1][10] = ready_o_1_10[0];
    data_o[1][11] = data_o_1_11[0];
    valid_o[1][11] = valid_o_1_11[0];
    ready_o[1][11] = ready_o_1_11[0];
    data_o[1][12] = data_o_1_12[0];
    valid_o[1][12] = valid_o_1_12[0];
    ready_o[1][12] = ready_o_1_12[0];
    data_o[1][13] = data_o_1_13[0];
    valid_o[1][13] = valid_o_1_13[0];
    ready_o[1][13] = ready_o_1_13[0];
    data_o[1][14] = data_o_1_14[0];
    valid_o[1][14] = valid_o_1_14[0];
    ready_o[1][14] = ready_o_1_14[0];
    data_o[1][15] = data_o_1_15[0];
    valid_o[1][15] = valid_o_1_15[0];
    ready_o[1][15] = ready_o_1_15[0];
    data_o[1][16] = data_o_1_16[0];
    valid_o[1][16] = valid_o_1_16[0];
    ready_o[1][16] = ready_o_1_16[0];
    data_o[1][17] = data_o_1_17[0];
    valid_o[1][17] = valid_o_1_17[0];
    ready_o[1][17] = ready_o_1_17[0];
    data_o[1][18] = data_o_1_18[0];
    valid_o[1][18] = valid_o_1_18[0];
    ready_o[1][18] = ready_o_1_18[0];
    data_o[1][19] = data_o_1_19[0];
    valid_o[1][19] = valid_o_1_19[0];
    ready_o[1][19] = ready_o_1_19[0];
    data_o[1][20] = data_o_1_20[0];
    valid_o[1][20] = valid_o_1_20[0];
    ready_o[1][20] = ready_o_1_20[0];
    data_o[1][21] = data_o_1_21[0];
    valid_o[1][21] = valid_o_1_21[0];
    ready_o[1][21] = ready_o_1_21[0];
    data_o[1][22] = data_o_1_22[0];
    valid_o[1][22] = valid_o_1_22[0];
    ready_o[1][22] = ready_o_1_22[0];
    data_o[1][23] = data_o_1_23[0];
    valid_o[1][23] = valid_o_1_23[0];
    ready_o[1][23] = ready_o_1_23[0];
    data_o[1][24] = data_o_1_24[0];
    valid_o[1][24] = valid_o_1_24[0];
    ready_o[1][24] = ready_o_1_24[0];
    data_o[2][0] = data_o_2_0[0];
    valid_o[2][0] = valid_o_2_0[0];
    ready_o[2][0] = ready_o_2_0[0];
    data_o[2][1] = data_o_2_1[0];
    valid_o[2][1] = valid_o_2_1[0];
    ready_o[2][1] = ready_o_2_1[0];
    data_o[2][2] = data_o_2_2[0];
    valid_o[2][2] = valid_o_2_2[0];
    ready_o[2][2] = ready_o_2_2[0];
    data_o[2][3] = data_o_2_3[0];
    valid_o[2][3] = valid_o_2_3[0];
    ready_o[2][3] = ready_o_2_3[0];
    data_o[2][4] = data_o_2_4[0];
    valid_o[2][4] = valid_o_2_4[0];
    ready_o[2][4] = ready_o_2_4[0];
    data_o[2][5] = data_o_2_5[0];
    valid_o[2][5] = valid_o_2_5[0];
    ready_o[2][5] = ready_o_2_5[0];
    data_o[2][6] = data_o_2_6[0];
    valid_o[2][6] = valid_o_2_6[0];
    ready_o[2][6] = ready_o_2_6[0];
    data_o[2][7] = data_o_2_7[0];
    valid_o[2][7] = valid_o_2_7[0];
    ready_o[2][7] = ready_o_2_7[0];
    data_o[2][8] = data_o_2_8[0];
    valid_o[2][8] = valid_o_2_8[0];
    ready_o[2][8] = ready_o_2_8[0];
    data_o[2][9] = data_o_2_9[0];
    valid_o[2][9] = valid_o_2_9[0];
    ready_o[2][9] = ready_o_2_9[0];
    data_o[2][10] = data_o_2_10[0];
    valid_o[2][10] = valid_o_2_10[0];
    ready_o[2][10] = ready_o_2_10[0];
    data_o[2][11] = data_o_2_11[0];
    valid_o[2][11] = valid_o_2_11[0];
    ready_o[2][11] = ready_o_2_11[0];
    data_o[2][12] = data_o_2_12[0];
    valid_o[2][12] = valid_o_2_12[0];
    ready_o[2][12] = ready_o_2_12[0];
    data_o[2][13] = data_o_2_13[0];
    valid_o[2][13] = valid_o_2_13[0];
    ready_o[2][13] = ready_o_2_13[0];
    data_o[2][14] = data_o_2_14[0];
    valid_o[2][14] = valid_o_2_14[0];
    ready_o[2][14] = ready_o_2_14[0];
    data_o[2][15] = data_o_2_15[0];
    valid_o[2][15] = valid_o_2_15[0];
    ready_o[2][15] = ready_o_2_15[0];
    data_o[2][16] = data_o_2_16[0];
    valid_o[2][16] = valid_o_2_16[0];
    ready_o[2][16] = ready_o_2_16[0];
    data_o[2][17] = data_o_2_17[0];
    valid_o[2][17] = valid_o_2_17[0];
    ready_o[2][17] = ready_o_2_17[0];
    data_o[2][18] = data_o_2_18[0];
    valid_o[2][18] = valid_o_2_18[0];
    ready_o[2][18] = ready_o_2_18[0];
    data_o[2][19] = data_o_2_19[0];
    valid_o[2][19] = valid_o_2_19[0];
    ready_o[2][19] = ready_o_2_19[0];
    data_o[2][20] = data_o_2_20[0];
    valid_o[2][20] = valid_o_2_20[0];
    ready_o[2][20] = ready_o_2_20[0];
    data_o[2][21] = data_o_2_21[0];
    valid_o[2][21] = valid_o_2_21[0];
    ready_o[2][21] = ready_o_2_21[0];
    data_o[2][22] = data_o_2_22[0];
    valid_o[2][22] = valid_o_2_22[0];
    ready_o[2][22] = ready_o_2_22[0];
    data_o[2][23] = data_o_2_23[0];
    valid_o[2][23] = valid_o_2_23[0];
    ready_o[2][23] = ready_o_2_23[0];
    data_o[2][24] = data_o_2_24[0];
    valid_o[2][24] = valid_o_2_24[0];
    ready_o[2][24] = ready_o_2_24[0];
    data_o[3][0] = data_o_3_0[0];
    valid_o[3][0] = valid_o_3_0[0];
    ready_o[3][0] = ready_o_3_0[0];
    data_o[3][1] = data_o_3_1[0];
    valid_o[3][1] = valid_o_3_1[0];
    ready_o[3][1] = ready_o_3_1[0];
    data_o[3][2] = data_o_3_2[0];
    valid_o[3][2] = valid_o_3_2[0];
    ready_o[3][2] = ready_o_3_2[0];
    data_o[3][3] = data_o_3_3[0];
    valid_o[3][3] = valid_o_3_3[0];
    ready_o[3][3] = ready_o_3_3[0];
    data_o[3][4] = data_o_3_4[0];
    valid_o[3][4] = valid_o_3_4[0];
    ready_o[3][4] = ready_o_3_4[0];
    data_o[3][5] = data_o_3_5[0];
    valid_o[3][5] = valid_o_3_5[0];
    ready_o[3][5] = ready_o_3_5[0];
    data_o[3][6] = data_o_3_6[0];
    valid_o[3][6] = valid_o_3_6[0];
    ready_o[3][6] = ready_o_3_6[0];
    data_o[3][7] = data_o_3_7[0];
    valid_o[3][7] = valid_o_3_7[0];
    ready_o[3][7] = ready_o_3_7[0];
    data_o[3][8] = data_o_3_8[0];
    valid_o[3][8] = valid_o_3_8[0];
    ready_o[3][8] = ready_o_3_8[0];
    data_o[3][9] = data_o_3_9[0];
    valid_o[3][9] = valid_o_3_9[0];
    ready_o[3][9] = ready_o_3_9[0];
    data_o[3][10] = data_o_3_10[0];
    valid_o[3][10] = valid_o_3_10[0];
    ready_o[3][10] = ready_o_3_10[0];
    data_o[3][11] = data_o_3_11[0];
    valid_o[3][11] = valid_o_3_11[0];
    ready_o[3][11] = ready_o_3_11[0];
    data_o[3][12] = data_o_3_12[0];
    valid_o[3][12] = valid_o_3_12[0];
    ready_o[3][12] = ready_o_3_12[0];
    data_o[3][13] = data_o_3_13[0];
    valid_o[3][13] = valid_o_3_13[0];
    ready_o[3][13] = ready_o_3_13[0];
    data_o[3][14] = data_o_3_14[0];
    valid_o[3][14] = valid_o_3_14[0];
    ready_o[3][14] = ready_o_3_14[0];
    data_o[3][15] = data_o_3_15[0];
    valid_o[3][15] = valid_o_3_15[0];
    ready_o[3][15] = ready_o_3_15[0];
    data_o[3][16] = data_o_3_16[0];
    valid_o[3][16] = valid_o_3_16[0];
    ready_o[3][16] = ready_o_3_16[0];
    data_o[3][17] = data_o_3_17[0];
    valid_o[3][17] = valid_o_3_17[0];
    ready_o[3][17] = ready_o_3_17[0];
    data_o[3][18] = data_o_3_18[0];
    valid_o[3][18] = valid_o_3_18[0];
    ready_o[3][18] = ready_o_3_18[0];
    data_o[3][19] = data_o_3_19[0];
    valid_o[3][19] = valid_o_3_19[0];
    ready_o[3][19] = ready_o_3_19[0];
    data_o[3][20] = data_o_3_20[0];
    valid_o[3][20] = valid_o_3_20[0];
    ready_o[3][20] = ready_o_3_20[0];
    data_o[3][21] = data_o_3_21[0];
    valid_o[3][21] = valid_o_3_21[0];
    ready_o[3][21] = ready_o_3_21[0];
    data_o[3][22] = data_o_3_22[0];
    valid_o[3][22] = valid_o_3_22[0];
    ready_o[3][22] = ready_o_3_22[0];
    data_o[3][23] = data_o_3_23[0];
    valid_o[3][23] = valid_o_3_23[0];
    ready_o[3][23] = ready_o_3_23[0];
    data_o[3][24] = data_o_3_24[0];
    valid_o[3][24] = valid_o_3_24[0];
    ready_o[3][24] = ready_o_3_24[0];
    data_o[4][0] = data_o_4_0[0];
    valid_o[4][0] = valid_o_4_0[0];
    ready_o[4][0] = ready_o_4_0[0];
    data_o[4][1] = data_o_4_1[0];
    valid_o[4][1] = valid_o_4_1[0];
    ready_o[4][1] = ready_o_4_1[0];
    data_o[4][2] = data_o_4_2[0];
    valid_o[4][2] = valid_o_4_2[0];
    ready_o[4][2] = ready_o_4_2[0];
    data_o[4][3] = data_o_4_3[0];
    valid_o[4][3] = valid_o_4_3[0];
    ready_o[4][3] = ready_o_4_3[0];
    data_o[4][4] = data_o_4_4[0];
    valid_o[4][4] = valid_o_4_4[0];
    ready_o[4][4] = ready_o_4_4[0];
    data_o[4][5] = data_o_4_5[0];
    valid_o[4][5] = valid_o_4_5[0];
    ready_o[4][5] = ready_o_4_5[0];
    data_o[4][6] = data_o_4_6[0];
    valid_o[4][6] = valid_o_4_6[0];
    ready_o[4][6] = ready_o_4_6[0];
    data_o[4][7] = data_o_4_7[0];
    valid_o[4][7] = valid_o_4_7[0];
    ready_o[4][7] = ready_o_4_7[0];
    data_o[4][8] = data_o_4_8[0];
    valid_o[4][8] = valid_o_4_8[0];
    ready_o[4][8] = ready_o_4_8[0];
    data_o[4][9] = data_o_4_9[0];
    valid_o[4][9] = valid_o_4_9[0];
    ready_o[4][9] = ready_o_4_9[0];
    data_o[4][10] = data_o_4_10[0];
    valid_o[4][10] = valid_o_4_10[0];
    ready_o[4][10] = ready_o_4_10[0];
    data_o[4][11] = data_o_4_11[0];
    valid_o[4][11] = valid_o_4_11[0];
    ready_o[4][11] = ready_o_4_11[0];
    data_o[4][12] = data_o_4_12[0];
    valid_o[4][12] = valid_o_4_12[0];
    ready_o[4][12] = ready_o_4_12[0];
    data_o[4][13] = data_o_4_13[0];
    valid_o[4][13] = valid_o_4_13[0];
    ready_o[4][13] = ready_o_4_13[0];
    data_o[4][14] = data_o_4_14[0];
    valid_o[4][14] = valid_o_4_14[0];
    ready_o[4][14] = ready_o_4_14[0];
    data_o[4][15] = data_o_4_15[0];
    valid_o[4][15] = valid_o_4_15[0];
    ready_o[4][15] = ready_o_4_15[0];
    data_o[4][16] = data_o_4_16[0];
    valid_o[4][16] = valid_o_4_16[0];
    ready_o[4][16] = ready_o_4_16[0];
    data_o[4][17] = data_o_4_17[0];
    valid_o[4][17] = valid_o_4_17[0];
    ready_o[4][17] = ready_o_4_17[0];
    data_o[4][18] = data_o_4_18[0];
    valid_o[4][18] = valid_o_4_18[0];
    ready_o[4][18] = ready_o_4_18[0];
    data_o[4][19] = data_o_4_19[0];
    valid_o[4][19] = valid_o_4_19[0];
    ready_o[4][19] = ready_o_4_19[0];
    data_o[4][20] = data_o_4_20[0];
    valid_o[4][20] = valid_o_4_20[0];
    ready_o[4][20] = ready_o_4_20[0];
    data_o[4][21] = data_o_4_21[0];
    valid_o[4][21] = valid_o_4_21[0];
    ready_o[4][21] = ready_o_4_21[0];
    data_o[4][22] = data_o_4_22[0];
    valid_o[4][22] = valid_o_4_22[0];
    ready_o[4][22] = ready_o_4_22[0];
    data_o[4][23] = data_o_4_23[0];
    valid_o[4][23] = valid_o_4_23[0];
    ready_o[4][23] = ready_o_4_23[0];
    data_o[4][24] = data_o_4_24[0];
    valid_o[4][24] = valid_o_4_24[0];
    ready_o[4][24] = ready_o_4_24[0];
    data_o[5][0] = data_o_5_0[0];
    valid_o[5][0] = valid_o_5_0[0];
    ready_o[5][0] = ready_o_5_0[0];
    data_o[5][1] = data_o_5_1[0];
    valid_o[5][1] = valid_o_5_1[0];
    ready_o[5][1] = ready_o_5_1[0];
    data_o[5][2] = data_o_5_2[0];
    valid_o[5][2] = valid_o_5_2[0];
    ready_o[5][2] = ready_o_5_2[0];
    data_o[5][3] = data_o_5_3[0];
    valid_o[5][3] = valid_o_5_3[0];
    ready_o[5][3] = ready_o_5_3[0];
    data_o[5][4] = data_o_5_4[0];
    valid_o[5][4] = valid_o_5_4[0];
    ready_o[5][4] = ready_o_5_4[0];
    data_o[5][5] = data_o_5_5[0];
    valid_o[5][5] = valid_o_5_5[0];
    ready_o[5][5] = ready_o_5_5[0];
    data_o[5][6] = data_o_5_6[0];
    valid_o[5][6] = valid_o_5_6[0];
    ready_o[5][6] = ready_o_5_6[0];
    data_o[5][7] = data_o_5_7[0];
    valid_o[5][7] = valid_o_5_7[0];
    ready_o[5][7] = ready_o_5_7[0];
    data_o[5][8] = data_o_5_8[0];
    valid_o[5][8] = valid_o_5_8[0];
    ready_o[5][8] = ready_o_5_8[0];
    data_o[5][9] = data_o_5_9[0];
    valid_o[5][9] = valid_o_5_9[0];
    ready_o[5][9] = ready_o_5_9[0];
    data_o[5][10] = data_o_5_10[0];
    valid_o[5][10] = valid_o_5_10[0];
    ready_o[5][10] = ready_o_5_10[0];
    data_o[5][11] = data_o_5_11[0];
    valid_o[5][11] = valid_o_5_11[0];
    ready_o[5][11] = ready_o_5_11[0];
    data_o[5][12] = data_o_5_12[0];
    valid_o[5][12] = valid_o_5_12[0];
    ready_o[5][12] = ready_o_5_12[0];
    data_o[5][13] = data_o_5_13[0];
    valid_o[5][13] = valid_o_5_13[0];
    ready_o[5][13] = ready_o_5_13[0];
    data_o[5][14] = data_o_5_14[0];
    valid_o[5][14] = valid_o_5_14[0];
    ready_o[5][14] = ready_o_5_14[0];
    data_o[5][15] = data_o_5_15[0];
    valid_o[5][15] = valid_o_5_15[0];
    ready_o[5][15] = ready_o_5_15[0];
    data_o[5][16] = data_o_5_16[0];
    valid_o[5][16] = valid_o_5_16[0];
    ready_o[5][16] = ready_o_5_16[0];
    data_o[5][17] = data_o_5_17[0];
    valid_o[5][17] = valid_o_5_17[0];
    ready_o[5][17] = ready_o_5_17[0];
    data_o[5][18] = data_o_5_18[0];
    valid_o[5][18] = valid_o_5_18[0];
    ready_o[5][18] = ready_o_5_18[0];
    data_o[5][19] = data_o_5_19[0];
    valid_o[5][19] = valid_o_5_19[0];
    ready_o[5][19] = ready_o_5_19[0];
    data_o[5][20] = data_o_5_20[0];
    valid_o[5][20] = valid_o_5_20[0];
    ready_o[5][20] = ready_o_5_20[0];
    data_o[5][21] = data_o_5_21[0];
    valid_o[5][21] = valid_o_5_21[0];
    ready_o[5][21] = ready_o_5_21[0];
    data_o[5][22] = data_o_5_22[0];
    valid_o[5][22] = valid_o_5_22[0];
    ready_o[5][22] = ready_o_5_22[0];
    data_o[5][23] = data_o_5_23[0];
    valid_o[5][23] = valid_o_5_23[0];
    ready_o[5][23] = ready_o_5_23[0];
    data_o[5][24] = data_o_5_24[0];
    valid_o[5][24] = valid_o_5_24[0];
    ready_o[5][24] = ready_o_5_24[0];
    data_o[6][0] = data_o_6_0[0];
    valid_o[6][0] = valid_o_6_0[0];
    ready_o[6][0] = ready_o_6_0[0];
    data_o[6][1] = data_o_6_1[0];
    valid_o[6][1] = valid_o_6_1[0];
    ready_o[6][1] = ready_o_6_1[0];
    data_o[6][2] = data_o_6_2[0];
    valid_o[6][2] = valid_o_6_2[0];
    ready_o[6][2] = ready_o_6_2[0];
    data_o[6][3] = data_o_6_3[0];
    valid_o[6][3] = valid_o_6_3[0];
    ready_o[6][3] = ready_o_6_3[0];
    data_o[6][4] = data_o_6_4[0];
    valid_o[6][4] = valid_o_6_4[0];
    ready_o[6][4] = ready_o_6_4[0];
    data_o[6][5] = data_o_6_5[0];
    valid_o[6][5] = valid_o_6_5[0];
    ready_o[6][5] = ready_o_6_5[0];
    data_o[6][6] = data_o_6_6[0];
    valid_o[6][6] = valid_o_6_6[0];
    ready_o[6][6] = ready_o_6_6[0];
    data_o[6][7] = data_o_6_7[0];
    valid_o[6][7] = valid_o_6_7[0];
    ready_o[6][7] = ready_o_6_7[0];
    data_o[6][8] = data_o_6_8[0];
    valid_o[6][8] = valid_o_6_8[0];
    ready_o[6][8] = ready_o_6_8[0];
    data_o[6][9] = data_o_6_9[0];
    valid_o[6][9] = valid_o_6_9[0];
    ready_o[6][9] = ready_o_6_9[0];
    data_o[6][10] = data_o_6_10[0];
    valid_o[6][10] = valid_o_6_10[0];
    ready_o[6][10] = ready_o_6_10[0];
    data_o[6][11] = data_o_6_11[0];
    valid_o[6][11] = valid_o_6_11[0];
    ready_o[6][11] = ready_o_6_11[0];
    data_o[6][12] = data_o_6_12[0];
    valid_o[6][12] = valid_o_6_12[0];
    ready_o[6][12] = ready_o_6_12[0];
    data_o[6][13] = data_o_6_13[0];
    valid_o[6][13] = valid_o_6_13[0];
    ready_o[6][13] = ready_o_6_13[0];
    data_o[6][14] = data_o_6_14[0];
    valid_o[6][14] = valid_o_6_14[0];
    ready_o[6][14] = ready_o_6_14[0];
    data_o[6][15] = data_o_6_15[0];
    valid_o[6][15] = valid_o_6_15[0];
    ready_o[6][15] = ready_o_6_15[0];
    data_o[6][16] = data_o_6_16[0];
    valid_o[6][16] = valid_o_6_16[0];
    ready_o[6][16] = ready_o_6_16[0];
    data_o[6][17] = data_o_6_17[0];
    valid_o[6][17] = valid_o_6_17[0];
    ready_o[6][17] = ready_o_6_17[0];
    data_o[6][18] = data_o_6_18[0];
    valid_o[6][18] = valid_o_6_18[0];
    ready_o[6][18] = ready_o_6_18[0];
    data_o[6][19] = data_o_6_19[0];
    valid_o[6][19] = valid_o_6_19[0];
    ready_o[6][19] = ready_o_6_19[0];
    data_o[6][20] = data_o_6_20[0];
    valid_o[6][20] = valid_o_6_20[0];
    ready_o[6][20] = ready_o_6_20[0];
    data_o[6][21] = data_o_6_21[0];
    valid_o[6][21] = valid_o_6_21[0];
    ready_o[6][21] = ready_o_6_21[0];
    data_o[6][22] = data_o_6_22[0];
    valid_o[6][22] = valid_o_6_22[0];
    ready_o[6][22] = ready_o_6_22[0];
    data_o[6][23] = data_o_6_23[0];
    valid_o[6][23] = valid_o_6_23[0];
    ready_o[6][23] = ready_o_6_23[0];
    data_o[6][24] = data_o_6_24[0];
    valid_o[6][24] = valid_o_6_24[0];
    ready_o[6][24] = ready_o_6_24[0];
    data_o[7][0] = data_o_7_0[0];
    valid_o[7][0] = valid_o_7_0[0];
    ready_o[7][0] = ready_o_7_0[0];
    data_o[7][1] = data_o_7_1[0];
    valid_o[7][1] = valid_o_7_1[0];
    ready_o[7][1] = ready_o_7_1[0];
    data_o[7][2] = data_o_7_2[0];
    valid_o[7][2] = valid_o_7_2[0];
    ready_o[7][2] = ready_o_7_2[0];
    data_o[7][3] = data_o_7_3[0];
    valid_o[7][3] = valid_o_7_3[0];
    ready_o[7][3] = ready_o_7_3[0];
    data_o[7][4] = data_o_7_4[0];
    valid_o[7][4] = valid_o_7_4[0];
    ready_o[7][4] = ready_o_7_4[0];
    data_o[7][5] = data_o_7_5[0];
    valid_o[7][5] = valid_o_7_5[0];
    ready_o[7][5] = ready_o_7_5[0];
    data_o[7][6] = data_o_7_6[0];
    valid_o[7][6] = valid_o_7_6[0];
    ready_o[7][6] = ready_o_7_6[0];
    data_o[7][7] = data_o_7_7[0];
    valid_o[7][7] = valid_o_7_7[0];
    ready_o[7][7] = ready_o_7_7[0];
    data_o[7][8] = data_o_7_8[0];
    valid_o[7][8] = valid_o_7_8[0];
    ready_o[7][8] = ready_o_7_8[0];
    data_o[7][9] = data_o_7_9[0];
    valid_o[7][9] = valid_o_7_9[0];
    ready_o[7][9] = ready_o_7_9[0];
    data_o[7][10] = data_o_7_10[0];
    valid_o[7][10] = valid_o_7_10[0];
    ready_o[7][10] = ready_o_7_10[0];
    data_o[7][11] = data_o_7_11[0];
    valid_o[7][11] = valid_o_7_11[0];
    ready_o[7][11] = ready_o_7_11[0];
    data_o[7][12] = data_o_7_12[0];
    valid_o[7][12] = valid_o_7_12[0];
    ready_o[7][12] = ready_o_7_12[0];
    data_o[7][13] = data_o_7_13[0];
    valid_o[7][13] = valid_o_7_13[0];
    ready_o[7][13] = ready_o_7_13[0];
    data_o[7][14] = data_o_7_14[0];
    valid_o[7][14] = valid_o_7_14[0];
    ready_o[7][14] = ready_o_7_14[0];
    data_o[7][15] = data_o_7_15[0];
    valid_o[7][15] = valid_o_7_15[0];
    ready_o[7][15] = ready_o_7_15[0];
    data_o[7][16] = data_o_7_16[0];
    valid_o[7][16] = valid_o_7_16[0];
    ready_o[7][16] = ready_o_7_16[0];
    data_o[7][17] = data_o_7_17[0];
    valid_o[7][17] = valid_o_7_17[0];
    ready_o[7][17] = ready_o_7_17[0];
    data_o[7][18] = data_o_7_18[0];
    valid_o[7][18] = valid_o_7_18[0];
    ready_o[7][18] = ready_o_7_18[0];
    data_o[7][19] = data_o_7_19[0];
    valid_o[7][19] = valid_o_7_19[0];
    ready_o[7][19] = ready_o_7_19[0];
    data_o[7][20] = data_o_7_20[0];
    valid_o[7][20] = valid_o_7_20[0];
    ready_o[7][20] = ready_o_7_20[0];
    data_o[7][21] = data_o_7_21[0];
    valid_o[7][21] = valid_o_7_21[0];
    ready_o[7][21] = ready_o_7_21[0];
    data_o[7][22] = data_o_7_22[0];
    valid_o[7][22] = valid_o_7_22[0];
    ready_o[7][22] = ready_o_7_22[0];
    data_o[7][23] = data_o_7_23[0];
    valid_o[7][23] = valid_o_7_23[0];
    ready_o[7][23] = ready_o_7_23[0];
    data_o[7][24] = data_o_7_24[0];
    valid_o[7][24] = valid_o_7_24[0];
    ready_o[7][24] = ready_o_7_24[0];
    data_o[8][0] = data_o_8_0[0];
    valid_o[8][0] = valid_o_8_0[0];
    ready_o[8][0] = ready_o_8_0[0];
    data_o[8][1] = data_o_8_1[0];
    valid_o[8][1] = valid_o_8_1[0];
    ready_o[8][1] = ready_o_8_1[0];
    data_o[8][2] = data_o_8_2[0];
    valid_o[8][2] = valid_o_8_2[0];
    ready_o[8][2] = ready_o_8_2[0];
    data_o[8][3] = data_o_8_3[0];
    valid_o[8][3] = valid_o_8_3[0];
    ready_o[8][3] = ready_o_8_3[0];
    data_o[8][4] = data_o_8_4[0];
    valid_o[8][4] = valid_o_8_4[0];
    ready_o[8][4] = ready_o_8_4[0];
    data_o[8][5] = data_o_8_5[0];
    valid_o[8][5] = valid_o_8_5[0];
    ready_o[8][5] = ready_o_8_5[0];
    data_o[8][6] = data_o_8_6[0];
    valid_o[8][6] = valid_o_8_6[0];
    ready_o[8][6] = ready_o_8_6[0];
    data_o[8][7] = data_o_8_7[0];
    valid_o[8][7] = valid_o_8_7[0];
    ready_o[8][7] = ready_o_8_7[0];
    data_o[8][8] = data_o_8_8[0];
    valid_o[8][8] = valid_o_8_8[0];
    ready_o[8][8] = ready_o_8_8[0];
    data_o[8][9] = data_o_8_9[0];
    valid_o[8][9] = valid_o_8_9[0];
    ready_o[8][9] = ready_o_8_9[0];
    data_o[8][10] = data_o_8_10[0];
    valid_o[8][10] = valid_o_8_10[0];
    ready_o[8][10] = ready_o_8_10[0];
    data_o[8][11] = data_o_8_11[0];
    valid_o[8][11] = valid_o_8_11[0];
    ready_o[8][11] = ready_o_8_11[0];
    data_o[8][12] = data_o_8_12[0];
    valid_o[8][12] = valid_o_8_12[0];
    ready_o[8][12] = ready_o_8_12[0];
    data_o[8][13] = data_o_8_13[0];
    valid_o[8][13] = valid_o_8_13[0];
    ready_o[8][13] = ready_o_8_13[0];
    data_o[8][14] = data_o_8_14[0];
    valid_o[8][14] = valid_o_8_14[0];
    ready_o[8][14] = ready_o_8_14[0];
    data_o[8][15] = data_o_8_15[0];
    valid_o[8][15] = valid_o_8_15[0];
    ready_o[8][15] = ready_o_8_15[0];
    data_o[8][16] = data_o_8_16[0];
    valid_o[8][16] = valid_o_8_16[0];
    ready_o[8][16] = ready_o_8_16[0];
    data_o[8][17] = data_o_8_17[0];
    valid_o[8][17] = valid_o_8_17[0];
    ready_o[8][17] = ready_o_8_17[0];
    data_o[8][18] = data_o_8_18[0];
    valid_o[8][18] = valid_o_8_18[0];
    ready_o[8][18] = ready_o_8_18[0];
    data_o[8][19] = data_o_8_19[0];
    valid_o[8][19] = valid_o_8_19[0];
    ready_o[8][19] = ready_o_8_19[0];
    data_o[8][20] = data_o_8_20[0];
    valid_o[8][20] = valid_o_8_20[0];
    ready_o[8][20] = ready_o_8_20[0];
    data_o[8][21] = data_o_8_21[0];
    valid_o[8][21] = valid_o_8_21[0];
    ready_o[8][21] = ready_o_8_21[0];
    data_o[8][22] = data_o_8_22[0];
    valid_o[8][22] = valid_o_8_22[0];
    ready_o[8][22] = ready_o_8_22[0];
    data_o[8][23] = data_o_8_23[0];
    valid_o[8][23] = valid_o_8_23[0];
    ready_o[8][23] = ready_o_8_23[0];
    data_o[8][24] = data_o_8_24[0];
    valid_o[8][24] = valid_o_8_24[0];
    ready_o[8][24] = ready_o_8_24[0];
    data_o[9][0] = data_o_9_0[0];
    valid_o[9][0] = valid_o_9_0[0];
    ready_o[9][0] = ready_o_9_0[0];
    data_o[9][1] = data_o_9_1[0];
    valid_o[9][1] = valid_o_9_1[0];
    ready_o[9][1] = ready_o_9_1[0];
    data_o[9][2] = data_o_9_2[0];
    valid_o[9][2] = valid_o_9_2[0];
    ready_o[9][2] = ready_o_9_2[0];
    data_o[9][3] = data_o_9_3[0];
    valid_o[9][3] = valid_o_9_3[0];
    ready_o[9][3] = ready_o_9_3[0];
    data_o[9][4] = data_o_9_4[0];
    valid_o[9][4] = valid_o_9_4[0];
    ready_o[9][4] = ready_o_9_4[0];
    data_o[9][5] = data_o_9_5[0];
    valid_o[9][5] = valid_o_9_5[0];
    ready_o[9][5] = ready_o_9_5[0];
    data_o[9][6] = data_o_9_6[0];
    valid_o[9][6] = valid_o_9_6[0];
    ready_o[9][6] = ready_o_9_6[0];
    data_o[9][7] = data_o_9_7[0];
    valid_o[9][7] = valid_o_9_7[0];
    ready_o[9][7] = ready_o_9_7[0];
    data_o[9][8] = data_o_9_8[0];
    valid_o[9][8] = valid_o_9_8[0];
    ready_o[9][8] = ready_o_9_8[0];
    data_o[9][9] = data_o_9_9[0];
    valid_o[9][9] = valid_o_9_9[0];
    ready_o[9][9] = ready_o_9_9[0];
    data_o[9][10] = data_o_9_10[0];
    valid_o[9][10] = valid_o_9_10[0];
    ready_o[9][10] = ready_o_9_10[0];
    data_o[9][11] = data_o_9_11[0];
    valid_o[9][11] = valid_o_9_11[0];
    ready_o[9][11] = ready_o_9_11[0];
    data_o[9][12] = data_o_9_12[0];
    valid_o[9][12] = valid_o_9_12[0];
    ready_o[9][12] = ready_o_9_12[0];
    data_o[9][13] = data_o_9_13[0];
    valid_o[9][13] = valid_o_9_13[0];
    ready_o[9][13] = ready_o_9_13[0];
    data_o[9][14] = data_o_9_14[0];
    valid_o[9][14] = valid_o_9_14[0];
    ready_o[9][14] = ready_o_9_14[0];
    data_o[9][15] = data_o_9_15[0];
    valid_o[9][15] = valid_o_9_15[0];
    ready_o[9][15] = ready_o_9_15[0];
    data_o[9][16] = data_o_9_16[0];
    valid_o[9][16] = valid_o_9_16[0];
    ready_o[9][16] = ready_o_9_16[0];
    data_o[9][17] = data_o_9_17[0];
    valid_o[9][17] = valid_o_9_17[0];
    ready_o[9][17] = ready_o_9_17[0];
    data_o[9][18] = data_o_9_18[0];
    valid_o[9][18] = valid_o_9_18[0];
    ready_o[9][18] = ready_o_9_18[0];
    data_o[9][19] = data_o_9_19[0];
    valid_o[9][19] = valid_o_9_19[0];
    ready_o[9][19] = ready_o_9_19[0];
    data_o[9][20] = data_o_9_20[0];
    valid_o[9][20] = valid_o_9_20[0];
    ready_o[9][20] = ready_o_9_20[0];
    data_o[9][21] = data_o_9_21[0];
    valid_o[9][21] = valid_o_9_21[0];
    ready_o[9][21] = ready_o_9_21[0];
    data_o[9][22] = data_o_9_22[0];
    valid_o[9][22] = valid_o_9_22[0];
    ready_o[9][22] = ready_o_9_22[0];
    data_o[9][23] = data_o_9_23[0];
    valid_o[9][23] = valid_o_9_23[0];
    ready_o[9][23] = ready_o_9_23[0];
    data_o[9][24] = data_o_9_24[0];
    valid_o[9][24] = valid_o_9_24[0];
    ready_o[9][24] = ready_o_9_24[0];
end

/*Router 0,0*/    
merge_router #(
    .input_mask                     (input_mask_0_0),
    .output_sel                     (output_sel_0_0)
)router0(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_0_0),
    .valid_i                        (valid_i_0_0),
    .ready_o                        (ready_o_0_0),
    .data_o                         (data_o_0_0),
    .valid_o                        (valid_o_0_0),
    .ready_i                        (ready_i_0_0)
);


always@(*) begin
    data_i_0_0[4] = data_o_0_1[3];
    valid_i_0_0[4] = valid_o_0_1[3];
    ready_i_0_0[4] = ready_o_0_1[3];
    data_i_0_0[2] = data_o_1_0[1];
    valid_i_0_0[2] = valid_o_1_0[1];
    ready_i_0_0[2] = ready_o_1_0[1];
    data_i_0_0[0] = data_i[0][0];
    valid_i_0_0[0] = valid_i[0][0];
    ready_i_0_0[0] = ready_i[0][0];
end


/*Router 0,1*/    
merge_router #(
    .input_mask                     (input_mask_0_1),
    .output_sel                     (output_sel_0_1)
)router10(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_0_1),
    .valid_i                        (valid_i_0_1),
    .ready_o                        (ready_o_0_1),
    .data_o                         (data_o_0_1),
    .valid_o                        (valid_o_0_1),
    .ready_i                        (ready_i_0_1)
);


always@(*) begin
    data_i_0_1[3] = data_o_0_0[4];
    valid_i_0_1[3] = valid_o_0_0[4];
    ready_i_0_1[3] = ready_o_0_0[4];
    data_i_0_1[4] = data_o_0_2[3];
    valid_i_0_1[4] = valid_o_0_2[3];
    ready_i_0_1[4] = ready_o_0_2[3];
    data_i_0_1[2] = data_o_1_1[1];
    valid_i_0_1[2] = valid_o_1_1[1];
    ready_i_0_1[2] = ready_o_1_1[1];
    data_i_0_1[0] = data_i[0][1];
    valid_i_0_1[0] = valid_i[0][1];
    ready_i_0_1[0] = ready_i[0][1];
end


/*Router 0,2*/    
merge_router #(
    .input_mask                     (input_mask_0_2),
    .output_sel                     (output_sel_0_2)
)router20(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_0_2),
    .valid_i                        (valid_i_0_2),
    .ready_o                        (ready_o_0_2),
    .data_o                         (data_o_0_2),
    .valid_o                        (valid_o_0_2),
    .ready_i                        (ready_i_0_2)
);


always@(*) begin
    data_i_0_2[3] = data_o_0_1[4];
    valid_i_0_2[3] = valid_o_0_1[4];
    ready_i_0_2[3] = ready_o_0_1[4];
    data_i_0_2[4] = data_o_0_3[3];
    valid_i_0_2[4] = valid_o_0_3[3];
    ready_i_0_2[4] = ready_o_0_3[3];
    data_i_0_2[2] = data_o_1_2[1];
    valid_i_0_2[2] = valid_o_1_2[1];
    ready_i_0_2[2] = ready_o_1_2[1];
    data_i_0_2[0] = data_i[0][2];
    valid_i_0_2[0] = valid_i[0][2];
    ready_i_0_2[0] = ready_i[0][2];
end


/*Router 0,3*/    
merge_router #(
    .input_mask                     (input_mask_0_3),
    .output_sel                     (output_sel_0_3)
)router30(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_0_3),
    .valid_i                        (valid_i_0_3),
    .ready_o                        (ready_o_0_3),
    .data_o                         (data_o_0_3),
    .valid_o                        (valid_o_0_3),
    .ready_i                        (ready_i_0_3)
);


always@(*) begin
    data_i_0_3[3] = data_o_0_2[4];
    valid_i_0_3[3] = valid_o_0_2[4];
    ready_i_0_3[3] = ready_o_0_2[4];
    data_i_0_3[4] = data_o_0_4[3];
    valid_i_0_3[4] = valid_o_0_4[3];
    ready_i_0_3[4] = ready_o_0_4[3];
    data_i_0_3[2] = data_o_1_3[1];
    valid_i_0_3[2] = valid_o_1_3[1];
    ready_i_0_3[2] = ready_o_1_3[1];
    data_i_0_3[0] = data_i[0][3];
    valid_i_0_3[0] = valid_i[0][3];
    ready_i_0_3[0] = ready_i[0][3];
end


/*Router 0,4*/    
merge_router #(
    .input_mask                     (input_mask_0_4),
    .output_sel                     (output_sel_0_4)
)router40(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_0_4),
    .valid_i                        (valid_i_0_4),
    .ready_o                        (ready_o_0_4),
    .data_o                         (data_o_0_4),
    .valid_o                        (valid_o_0_4),
    .ready_i                        (ready_i_0_4)
);


always@(*) begin
    data_i_0_4[3] = data_o_0_3[4];
    valid_i_0_4[3] = valid_o_0_3[4];
    ready_i_0_4[3] = ready_o_0_3[4];
    data_i_0_4[4] = data_o_0_5[3];
    valid_i_0_4[4] = valid_o_0_5[3];
    ready_i_0_4[4] = ready_o_0_5[3];
    data_i_0_4[2] = data_o_1_4[1];
    valid_i_0_4[2] = valid_o_1_4[1];
    ready_i_0_4[2] = ready_o_1_4[1];
    data_i_0_4[0] = data_i[0][4];
    valid_i_0_4[0] = valid_i[0][4];
    ready_i_0_4[0] = ready_i[0][4];
end


/*Router 0,5*/    
merge_router #(
    .input_mask                     (input_mask_0_5),
    .output_sel                     (output_sel_0_5)
)router50(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_0_5),
    .valid_i                        (valid_i_0_5),
    .ready_o                        (ready_o_0_5),
    .data_o                         (data_o_0_5),
    .valid_o                        (valid_o_0_5),
    .ready_i                        (ready_i_0_5)
);


always@(*) begin
    data_i_0_5[3] = data_o_0_4[4];
    valid_i_0_5[3] = valid_o_0_4[4];
    ready_i_0_5[3] = ready_o_0_4[4];
    data_i_0_5[4] = data_o_0_6[3];
    valid_i_0_5[4] = valid_o_0_6[3];
    ready_i_0_5[4] = ready_o_0_6[3];
    data_i_0_5[2] = data_o_1_5[1];
    valid_i_0_5[2] = valid_o_1_5[1];
    ready_i_0_5[2] = ready_o_1_5[1];
    data_i_0_5[0] = data_i[0][5];
    valid_i_0_5[0] = valid_i[0][5];
    ready_i_0_5[0] = ready_i[0][5];
end


/*Router 0,6*/    
merge_router #(
    .input_mask                     (input_mask_0_6),
    .output_sel                     (output_sel_0_6)
)router60(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_0_6),
    .valid_i                        (valid_i_0_6),
    .ready_o                        (ready_o_0_6),
    .data_o                         (data_o_0_6),
    .valid_o                        (valid_o_0_6),
    .ready_i                        (ready_i_0_6)
);


always@(*) begin
    data_i_0_6[3] = data_o_0_5[4];
    valid_i_0_6[3] = valid_o_0_5[4];
    ready_i_0_6[3] = ready_o_0_5[4];
    data_i_0_6[4] = data_o_0_7[3];
    valid_i_0_6[4] = valid_o_0_7[3];
    ready_i_0_6[4] = ready_o_0_7[3];
    data_i_0_6[2] = data_o_1_6[1];
    valid_i_0_6[2] = valid_o_1_6[1];
    ready_i_0_6[2] = ready_o_1_6[1];
    data_i_0_6[0] = data_i[0][6];
    valid_i_0_6[0] = valid_i[0][6];
    ready_i_0_6[0] = ready_i[0][6];
end


/*Router 0,7*/    
merge_router #(
    .input_mask                     (input_mask_0_7),
    .output_sel                     (output_sel_0_7)
)router70(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_0_7),
    .valid_i                        (valid_i_0_7),
    .ready_o                        (ready_o_0_7),
    .data_o                         (data_o_0_7),
    .valid_o                        (valid_o_0_7),
    .ready_i                        (ready_i_0_7)
);


always@(*) begin
    data_i_0_7[3] = data_o_0_6[4];
    valid_i_0_7[3] = valid_o_0_6[4];
    ready_i_0_7[3] = ready_o_0_6[4];
    data_i_0_7[4] = data_o_0_8[3];
    valid_i_0_7[4] = valid_o_0_8[3];
    ready_i_0_7[4] = ready_o_0_8[3];
    data_i_0_7[2] = data_o_1_7[1];
    valid_i_0_7[2] = valid_o_1_7[1];
    ready_i_0_7[2] = ready_o_1_7[1];
    data_i_0_7[0] = data_i[0][7];
    valid_i_0_7[0] = valid_i[0][7];
    ready_i_0_7[0] = ready_i[0][7];
end


/*Router 0,8*/    
merge_router #(
    .input_mask                     (input_mask_0_8),
    .output_sel                     (output_sel_0_8)
)router80(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_0_8),
    .valid_i                        (valid_i_0_8),
    .ready_o                        (ready_o_0_8),
    .data_o                         (data_o_0_8),
    .valid_o                        (valid_o_0_8),
    .ready_i                        (ready_i_0_8)
);


always@(*) begin
    data_i_0_8[3] = data_o_0_7[4];
    valid_i_0_8[3] = valid_o_0_7[4];
    ready_i_0_8[3] = ready_o_0_7[4];
    data_i_0_8[4] = data_o_0_9[3];
    valid_i_0_8[4] = valid_o_0_9[3];
    ready_i_0_8[4] = ready_o_0_9[3];
    data_i_0_8[2] = data_o_1_8[1];
    valid_i_0_8[2] = valid_o_1_8[1];
    ready_i_0_8[2] = ready_o_1_8[1];
    data_i_0_8[0] = data_i[0][8];
    valid_i_0_8[0] = valid_i[0][8];
    ready_i_0_8[0] = ready_i[0][8];
end


/*Router 0,9*/    
merge_router #(
    .input_mask                     (input_mask_0_9),
    .output_sel                     (output_sel_0_9)
)router90(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_0_9),
    .valid_i                        (valid_i_0_9),
    .ready_o                        (ready_o_0_9),
    .data_o                         (data_o_0_9),
    .valid_o                        (valid_o_0_9),
    .ready_i                        (ready_i_0_9)
);


always@(*) begin
    data_i_0_9[3] = data_o_0_8[4];
    valid_i_0_9[3] = valid_o_0_8[4];
    ready_i_0_9[3] = ready_o_0_8[4];
    data_i_0_9[4] = data_o_0_10[3];
    valid_i_0_9[4] = valid_o_0_10[3];
    ready_i_0_9[4] = ready_o_0_10[3];
    data_i_0_9[2] = data_o_1_9[1];
    valid_i_0_9[2] = valid_o_1_9[1];
    ready_i_0_9[2] = ready_o_1_9[1];
    data_i_0_9[0] = data_i[0][9];
    valid_i_0_9[0] = valid_i[0][9];
    ready_i_0_9[0] = ready_i[0][9];
end


/*Router 0,10*/    
merge_router #(
    .input_mask                     (input_mask_0_10),
    .output_sel                     (output_sel_0_10)
)router100(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_0_10),
    .valid_i                        (valid_i_0_10),
    .ready_o                        (ready_o_0_10),
    .data_o                         (data_o_0_10),
    .valid_o                        (valid_o_0_10),
    .ready_i                        (ready_i_0_10)
);


always@(*) begin
    data_i_0_10[3] = data_o_0_9[4];
    valid_i_0_10[3] = valid_o_0_9[4];
    ready_i_0_10[3] = ready_o_0_9[4];
    data_i_0_10[4] = data_o_0_11[3];
    valid_i_0_10[4] = valid_o_0_11[3];
    ready_i_0_10[4] = ready_o_0_11[3];
    data_i_0_10[2] = data_o_1_10[1];
    valid_i_0_10[2] = valid_o_1_10[1];
    ready_i_0_10[2] = ready_o_1_10[1];
    data_i_0_10[0] = data_i[0][10];
    valid_i_0_10[0] = valid_i[0][10];
    ready_i_0_10[0] = ready_i[0][10];
end


/*Router 0,11*/    
merge_router #(
    .input_mask                     (input_mask_0_11),
    .output_sel                     (output_sel_0_11)
)router110(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_0_11),
    .valid_i                        (valid_i_0_11),
    .ready_o                        (ready_o_0_11),
    .data_o                         (data_o_0_11),
    .valid_o                        (valid_o_0_11),
    .ready_i                        (ready_i_0_11)
);


always@(*) begin
    data_i_0_11[3] = data_o_0_10[4];
    valid_i_0_11[3] = valid_o_0_10[4];
    ready_i_0_11[3] = ready_o_0_10[4];
    data_i_0_11[4] = data_o_0_12[3];
    valid_i_0_11[4] = valid_o_0_12[3];
    ready_i_0_11[4] = ready_o_0_12[3];
    data_i_0_11[2] = data_o_1_11[1];
    valid_i_0_11[2] = valid_o_1_11[1];
    ready_i_0_11[2] = ready_o_1_11[1];
    data_i_0_11[0] = data_i[0][11];
    valid_i_0_11[0] = valid_i[0][11];
    ready_i_0_11[0] = ready_i[0][11];
end


/*Router 0,12*/    
merge_router #(
    .input_mask                     (input_mask_0_12),
    .output_sel                     (output_sel_0_12)
)router120(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_0_12),
    .valid_i                        (valid_i_0_12),
    .ready_o                        (ready_o_0_12),
    .data_o                         (data_o_0_12),
    .valid_o                        (valid_o_0_12),
    .ready_i                        (ready_i_0_12)
);


always@(*) begin
    data_i_0_12[3] = data_o_0_11[4];
    valid_i_0_12[3] = valid_o_0_11[4];
    ready_i_0_12[3] = ready_o_0_11[4];
    data_i_0_12[4] = data_o_0_13[3];
    valid_i_0_12[4] = valid_o_0_13[3];
    ready_i_0_12[4] = ready_o_0_13[3];
    data_i_0_12[2] = data_o_1_12[1];
    valid_i_0_12[2] = valid_o_1_12[1];
    ready_i_0_12[2] = ready_o_1_12[1];
    data_i_0_12[0] = data_i[0][12];
    valid_i_0_12[0] = valid_i[0][12];
    ready_i_0_12[0] = ready_i[0][12];
end


/*Router 0,13*/    
merge_router #(
    .input_mask                     (input_mask_0_13),
    .output_sel                     (output_sel_0_13)
)router130(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_0_13),
    .valid_i                        (valid_i_0_13),
    .ready_o                        (ready_o_0_13),
    .data_o                         (data_o_0_13),
    .valid_o                        (valid_o_0_13),
    .ready_i                        (ready_i_0_13)
);


always@(*) begin
    data_i_0_13[3] = data_o_0_12[4];
    valid_i_0_13[3] = valid_o_0_12[4];
    ready_i_0_13[3] = ready_o_0_12[4];
    data_i_0_13[4] = data_o_0_14[3];
    valid_i_0_13[4] = valid_o_0_14[3];
    ready_i_0_13[4] = ready_o_0_14[3];
    data_i_0_13[2] = data_o_1_13[1];
    valid_i_0_13[2] = valid_o_1_13[1];
    ready_i_0_13[2] = ready_o_1_13[1];
    data_i_0_13[0] = data_i[0][13];
    valid_i_0_13[0] = valid_i[0][13];
    ready_i_0_13[0] = ready_i[0][13];
end


/*Router 0,14*/    
merge_router #(
    .input_mask                     (input_mask_0_14),
    .output_sel                     (output_sel_0_14)
)router140(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_0_14),
    .valid_i                        (valid_i_0_14),
    .ready_o                        (ready_o_0_14),
    .data_o                         (data_o_0_14),
    .valid_o                        (valid_o_0_14),
    .ready_i                        (ready_i_0_14)
);


always@(*) begin
    data_i_0_14[3] = data_o_0_13[4];
    valid_i_0_14[3] = valid_o_0_13[4];
    ready_i_0_14[3] = ready_o_0_13[4];
    data_i_0_14[4] = data_o_0_15[3];
    valid_i_0_14[4] = valid_o_0_15[3];
    ready_i_0_14[4] = ready_o_0_15[3];
    data_i_0_14[2] = data_o_1_14[1];
    valid_i_0_14[2] = valid_o_1_14[1];
    ready_i_0_14[2] = ready_o_1_14[1];
    data_i_0_14[0] = data_i[0][14];
    valid_i_0_14[0] = valid_i[0][14];
    ready_i_0_14[0] = ready_i[0][14];
end


/*Router 0,15*/    
merge_router #(
    .input_mask                     (input_mask_0_15),
    .output_sel                     (output_sel_0_15)
)router150(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_0_15),
    .valid_i                        (valid_i_0_15),
    .ready_o                        (ready_o_0_15),
    .data_o                         (data_o_0_15),
    .valid_o                        (valid_o_0_15),
    .ready_i                        (ready_i_0_15)
);


always@(*) begin
    data_i_0_15[3] = data_o_0_14[4];
    valid_i_0_15[3] = valid_o_0_14[4];
    ready_i_0_15[3] = ready_o_0_14[4];
    data_i_0_15[4] = data_o_0_16[3];
    valid_i_0_15[4] = valid_o_0_16[3];
    ready_i_0_15[4] = ready_o_0_16[3];
    data_i_0_15[2] = data_o_1_15[1];
    valid_i_0_15[2] = valid_o_1_15[1];
    ready_i_0_15[2] = ready_o_1_15[1];
    data_i_0_15[0] = data_i[0][15];
    valid_i_0_15[0] = valid_i[0][15];
    ready_i_0_15[0] = ready_i[0][15];
end


/*Router 0,16*/    
merge_router #(
    .input_mask                     (input_mask_0_16),
    .output_sel                     (output_sel_0_16)
)router160(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_0_16),
    .valid_i                        (valid_i_0_16),
    .ready_o                        (ready_o_0_16),
    .data_o                         (data_o_0_16),
    .valid_o                        (valid_o_0_16),
    .ready_i                        (ready_i_0_16)
);


always@(*) begin
    data_i_0_16[3] = data_o_0_15[4];
    valid_i_0_16[3] = valid_o_0_15[4];
    ready_i_0_16[3] = ready_o_0_15[4];
    data_i_0_16[4] = data_o_0_17[3];
    valid_i_0_16[4] = valid_o_0_17[3];
    ready_i_0_16[4] = ready_o_0_17[3];
    data_i_0_16[2] = data_o_1_16[1];
    valid_i_0_16[2] = valid_o_1_16[1];
    ready_i_0_16[2] = ready_o_1_16[1];
    data_i_0_16[0] = data_i[0][16];
    valid_i_0_16[0] = valid_i[0][16];
    ready_i_0_16[0] = ready_i[0][16];
end


/*Router 0,17*/    
merge_router #(
    .input_mask                     (input_mask_0_17),
    .output_sel                     (output_sel_0_17)
)router170(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_0_17),
    .valid_i                        (valid_i_0_17),
    .ready_o                        (ready_o_0_17),
    .data_o                         (data_o_0_17),
    .valid_o                        (valid_o_0_17),
    .ready_i                        (ready_i_0_17)
);


always@(*) begin
    data_i_0_17[3] = data_o_0_16[4];
    valid_i_0_17[3] = valid_o_0_16[4];
    ready_i_0_17[3] = ready_o_0_16[4];
    data_i_0_17[4] = data_o_0_18[3];
    valid_i_0_17[4] = valid_o_0_18[3];
    ready_i_0_17[4] = ready_o_0_18[3];
    data_i_0_17[2] = data_o_1_17[1];
    valid_i_0_17[2] = valid_o_1_17[1];
    ready_i_0_17[2] = ready_o_1_17[1];
    data_i_0_17[0] = data_i[0][17];
    valid_i_0_17[0] = valid_i[0][17];
    ready_i_0_17[0] = ready_i[0][17];
end


/*Router 0,18*/    
merge_router #(
    .input_mask                     (input_mask_0_18),
    .output_sel                     (output_sel_0_18)
)router180(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_0_18),
    .valid_i                        (valid_i_0_18),
    .ready_o                        (ready_o_0_18),
    .data_o                         (data_o_0_18),
    .valid_o                        (valid_o_0_18),
    .ready_i                        (ready_i_0_18)
);


always@(*) begin
    data_i_0_18[3] = data_o_0_17[4];
    valid_i_0_18[3] = valid_o_0_17[4];
    ready_i_0_18[3] = ready_o_0_17[4];
    data_i_0_18[4] = data_o_0_19[3];
    valid_i_0_18[4] = valid_o_0_19[3];
    ready_i_0_18[4] = ready_o_0_19[3];
    data_i_0_18[2] = data_o_1_18[1];
    valid_i_0_18[2] = valid_o_1_18[1];
    ready_i_0_18[2] = ready_o_1_18[1];
    data_i_0_18[0] = data_i[0][18];
    valid_i_0_18[0] = valid_i[0][18];
    ready_i_0_18[0] = ready_i[0][18];
end


/*Router 0,19*/    
merge_router #(
    .input_mask                     (input_mask_0_19),
    .output_sel                     (output_sel_0_19)
)router190(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_0_19),
    .valid_i                        (valid_i_0_19),
    .ready_o                        (ready_o_0_19),
    .data_o                         (data_o_0_19),
    .valid_o                        (valid_o_0_19),
    .ready_i                        (ready_i_0_19)
);


always@(*) begin
    data_i_0_19[3] = data_o_0_18[4];
    valid_i_0_19[3] = valid_o_0_18[4];
    ready_i_0_19[3] = ready_o_0_18[4];
    data_i_0_19[4] = data_o_0_20[3];
    valid_i_0_19[4] = valid_o_0_20[3];
    ready_i_0_19[4] = ready_o_0_20[3];
    data_i_0_19[2] = data_o_1_19[1];
    valid_i_0_19[2] = valid_o_1_19[1];
    ready_i_0_19[2] = ready_o_1_19[1];
    data_i_0_19[0] = data_i[0][19];
    valid_i_0_19[0] = valid_i[0][19];
    ready_i_0_19[0] = ready_i[0][19];
end


/*Router 0,20*/    
merge_router #(
    .input_mask                     (input_mask_0_20),
    .output_sel                     (output_sel_0_20)
)router200(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_0_20),
    .valid_i                        (valid_i_0_20),
    .ready_o                        (ready_o_0_20),
    .data_o                         (data_o_0_20),
    .valid_o                        (valid_o_0_20),
    .ready_i                        (ready_i_0_20)
);


always@(*) begin
    data_i_0_20[3] = data_o_0_19[4];
    valid_i_0_20[3] = valid_o_0_19[4];
    ready_i_0_20[3] = ready_o_0_19[4];
    data_i_0_20[4] = data_o_0_21[3];
    valid_i_0_20[4] = valid_o_0_21[3];
    ready_i_0_20[4] = ready_o_0_21[3];
    data_i_0_20[2] = data_o_1_20[1];
    valid_i_0_20[2] = valid_o_1_20[1];
    ready_i_0_20[2] = ready_o_1_20[1];
    data_i_0_20[0] = data_i[0][20];
    valid_i_0_20[0] = valid_i[0][20];
    ready_i_0_20[0] = ready_i[0][20];
end


/*Router 0,21*/    
merge_router #(
    .input_mask                     (input_mask_0_21),
    .output_sel                     (output_sel_0_21)
)router210(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_0_21),
    .valid_i                        (valid_i_0_21),
    .ready_o                        (ready_o_0_21),
    .data_o                         (data_o_0_21),
    .valid_o                        (valid_o_0_21),
    .ready_i                        (ready_i_0_21)
);


always@(*) begin
    data_i_0_21[3] = data_o_0_20[4];
    valid_i_0_21[3] = valid_o_0_20[4];
    ready_i_0_21[3] = ready_o_0_20[4];
    data_i_0_21[4] = data_o_0_22[3];
    valid_i_0_21[4] = valid_o_0_22[3];
    ready_i_0_21[4] = ready_o_0_22[3];
    data_i_0_21[2] = data_o_1_21[1];
    valid_i_0_21[2] = valid_o_1_21[1];
    ready_i_0_21[2] = ready_o_1_21[1];
    data_i_0_21[0] = data_i[0][21];
    valid_i_0_21[0] = valid_i[0][21];
    ready_i_0_21[0] = ready_i[0][21];
end


/*Router 0,22*/    
merge_router #(
    .input_mask                     (input_mask_0_22),
    .output_sel                     (output_sel_0_22)
)router220(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_0_22),
    .valid_i                        (valid_i_0_22),
    .ready_o                        (ready_o_0_22),
    .data_o                         (data_o_0_22),
    .valid_o                        (valid_o_0_22),
    .ready_i                        (ready_i_0_22)
);


always@(*) begin
    data_i_0_22[3] = data_o_0_21[4];
    valid_i_0_22[3] = valid_o_0_21[4];
    ready_i_0_22[3] = ready_o_0_21[4];
    data_i_0_22[4] = data_o_0_23[3];
    valid_i_0_22[4] = valid_o_0_23[3];
    ready_i_0_22[4] = ready_o_0_23[3];
    data_i_0_22[2] = data_o_1_22[1];
    valid_i_0_22[2] = valid_o_1_22[1];
    ready_i_0_22[2] = ready_o_1_22[1];
    data_i_0_22[0] = data_i[0][22];
    valid_i_0_22[0] = valid_i[0][22];
    ready_i_0_22[0] = ready_i[0][22];
end


/*Router 0,23*/    
merge_router #(
    .input_mask                     (input_mask_0_23),
    .output_sel                     (output_sel_0_23)
)router230(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_0_23),
    .valid_i                        (valid_i_0_23),
    .ready_o                        (ready_o_0_23),
    .data_o                         (data_o_0_23),
    .valid_o                        (valid_o_0_23),
    .ready_i                        (ready_i_0_23)
);


always@(*) begin
    data_i_0_23[3] = data_o_0_22[4];
    valid_i_0_23[3] = valid_o_0_22[4];
    ready_i_0_23[3] = ready_o_0_22[4];
    data_i_0_23[4] = data_o_0_24[3];
    valid_i_0_23[4] = valid_o_0_24[3];
    ready_i_0_23[4] = ready_o_0_24[3];
    data_i_0_23[2] = data_o_1_23[1];
    valid_i_0_23[2] = valid_o_1_23[1];
    ready_i_0_23[2] = ready_o_1_23[1];
    data_i_0_23[0] = data_i[0][23];
    valid_i_0_23[0] = valid_i[0][23];
    ready_i_0_23[0] = ready_i[0][23];
end


/*Router 0,24*/    
merge_router #(
    .input_mask                     (input_mask_0_24),
    .output_sel                     (output_sel_0_24)
)router240(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_0_24),
    .valid_i                        (valid_i_0_24),
    .ready_o                        (ready_o_0_24),
    .data_o                         (data_o_0_24),
    .valid_o                        (valid_o_0_24),
    .ready_i                        (ready_i_0_24)
);


always@(*) begin
    data_i_0_24[3] = data_o_0_23[4];
    valid_i_0_24[3] = valid_o_0_23[4];
    ready_i_0_24[3] = ready_o_0_23[4];
    data_i_0_24[2] = data_o_1_24[1];
    valid_i_0_24[2] = valid_o_1_24[1];
    ready_i_0_24[2] = ready_o_1_24[1];
    data_i_0_24[0] = data_i[0][24];
    valid_i_0_24[0] = valid_i[0][24];
    ready_i_0_24[0] = ready_i[0][24];
end


/*Router 1,0*/    
merge_router #(
    .input_mask                     (input_mask_1_0),
    .output_sel                     (output_sel_1_0)
)router1(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_1_0),
    .valid_i                        (valid_i_1_0),
    .ready_o                        (ready_o_1_0),
    .data_o                         (data_o_1_0),
    .valid_o                        (valid_o_1_0),
    .ready_i                        (ready_i_1_0)
);


always@(*) begin
    data_i_1_0[4] = data_o_1_1[3];
    valid_i_1_0[4] = valid_o_1_1[3];
    ready_i_1_0[4] = ready_o_1_1[3];
    data_i_1_0[1] = data_o_0_0[2];
    valid_i_1_0[1] = valid_o_0_0[2];
    ready_i_1_0[1] = ready_o_0_0[2];
    data_i_1_0[2] = data_o_2_0[1];
    valid_i_1_0[2] = valid_o_2_0[1];
    ready_i_1_0[2] = ready_o_2_0[1];
    data_i_1_0[0] = data_i[1][0];
    valid_i_1_0[0] = valid_i[1][0];
    ready_i_1_0[0] = ready_i[1][0];
end


/*Router 1,1*/    
merge_router #(
    .input_mask                     (input_mask_1_1),
    .output_sel                     (output_sel_1_1)
)router11(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_1_1),
    .valid_i                        (valid_i_1_1),
    .ready_o                        (ready_o_1_1),
    .data_o                         (data_o_1_1),
    .valid_o                        (valid_o_1_1),
    .ready_i                        (ready_i_1_1)
);


always@(*) begin
    data_i_1_1[3] = data_o_1_0[4];
    valid_i_1_1[3] = valid_o_1_0[4];
    ready_i_1_1[3] = ready_o_1_0[4];
    data_i_1_1[4] = data_o_1_2[3];
    valid_i_1_1[4] = valid_o_1_2[3];
    ready_i_1_1[4] = ready_o_1_2[3];
    data_i_1_1[1] = data_o_0_1[2];
    valid_i_1_1[1] = valid_o_0_1[2];
    ready_i_1_1[1] = ready_o_0_1[2];
    data_i_1_1[2] = data_o_2_1[1];
    valid_i_1_1[2] = valid_o_2_1[1];
    ready_i_1_1[2] = ready_o_2_1[1];
    data_i_1_1[0] = data_i[1][1];
    valid_i_1_1[0] = valid_i[1][1];
    ready_i_1_1[0] = ready_i[1][1];
end


/*Router 1,2*/    
merge_router #(
    .input_mask                     (input_mask_1_2),
    .output_sel                     (output_sel_1_2)
)router21(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_1_2),
    .valid_i                        (valid_i_1_2),
    .ready_o                        (ready_o_1_2),
    .data_o                         (data_o_1_2),
    .valid_o                        (valid_o_1_2),
    .ready_i                        (ready_i_1_2)
);


always@(*) begin
    data_i_1_2[3] = data_o_1_1[4];
    valid_i_1_2[3] = valid_o_1_1[4];
    ready_i_1_2[3] = ready_o_1_1[4];
    data_i_1_2[4] = data_o_1_3[3];
    valid_i_1_2[4] = valid_o_1_3[3];
    ready_i_1_2[4] = ready_o_1_3[3];
    data_i_1_2[1] = data_o_0_2[2];
    valid_i_1_2[1] = valid_o_0_2[2];
    ready_i_1_2[1] = ready_o_0_2[2];
    data_i_1_2[2] = data_o_2_2[1];
    valid_i_1_2[2] = valid_o_2_2[1];
    ready_i_1_2[2] = ready_o_2_2[1];
    data_i_1_2[0] = data_i[1][2];
    valid_i_1_2[0] = valid_i[1][2];
    ready_i_1_2[0] = ready_i[1][2];
end


/*Router 1,3*/    
merge_router #(
    .input_mask                     (input_mask_1_3),
    .output_sel                     (output_sel_1_3)
)router31(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_1_3),
    .valid_i                        (valid_i_1_3),
    .ready_o                        (ready_o_1_3),
    .data_o                         (data_o_1_3),
    .valid_o                        (valid_o_1_3),
    .ready_i                        (ready_i_1_3)
);


always@(*) begin
    data_i_1_3[3] = data_o_1_2[4];
    valid_i_1_3[3] = valid_o_1_2[4];
    ready_i_1_3[3] = ready_o_1_2[4];
    data_i_1_3[4] = data_o_1_4[3];
    valid_i_1_3[4] = valid_o_1_4[3];
    ready_i_1_3[4] = ready_o_1_4[3];
    data_i_1_3[1] = data_o_0_3[2];
    valid_i_1_3[1] = valid_o_0_3[2];
    ready_i_1_3[1] = ready_o_0_3[2];
    data_i_1_3[2] = data_o_2_3[1];
    valid_i_1_3[2] = valid_o_2_3[1];
    ready_i_1_3[2] = ready_o_2_3[1];
    data_i_1_3[0] = data_i[1][3];
    valid_i_1_3[0] = valid_i[1][3];
    ready_i_1_3[0] = ready_i[1][3];
end


/*Router 1,4*/    
merge_router #(
    .input_mask                     (input_mask_1_4),
    .output_sel                     (output_sel_1_4)
)router41(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_1_4),
    .valid_i                        (valid_i_1_4),
    .ready_o                        (ready_o_1_4),
    .data_o                         (data_o_1_4),
    .valid_o                        (valid_o_1_4),
    .ready_i                        (ready_i_1_4)
);


always@(*) begin
    data_i_1_4[3] = data_o_1_3[4];
    valid_i_1_4[3] = valid_o_1_3[4];
    ready_i_1_4[3] = ready_o_1_3[4];
    data_i_1_4[4] = data_o_1_5[3];
    valid_i_1_4[4] = valid_o_1_5[3];
    ready_i_1_4[4] = ready_o_1_5[3];
    data_i_1_4[1] = data_o_0_4[2];
    valid_i_1_4[1] = valid_o_0_4[2];
    ready_i_1_4[1] = ready_o_0_4[2];
    data_i_1_4[2] = data_o_2_4[1];
    valid_i_1_4[2] = valid_o_2_4[1];
    ready_i_1_4[2] = ready_o_2_4[1];
    data_i_1_4[0] = data_i[1][4];
    valid_i_1_4[0] = valid_i[1][4];
    ready_i_1_4[0] = ready_i[1][4];
end


/*Router 1,5*/    
merge_router #(
    .input_mask                     (input_mask_1_5),
    .output_sel                     (output_sel_1_5)
)router51(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_1_5),
    .valid_i                        (valid_i_1_5),
    .ready_o                        (ready_o_1_5),
    .data_o                         (data_o_1_5),
    .valid_o                        (valid_o_1_5),
    .ready_i                        (ready_i_1_5)
);


always@(*) begin
    data_i_1_5[3] = data_o_1_4[4];
    valid_i_1_5[3] = valid_o_1_4[4];
    ready_i_1_5[3] = ready_o_1_4[4];
    data_i_1_5[4] = data_o_1_6[3];
    valid_i_1_5[4] = valid_o_1_6[3];
    ready_i_1_5[4] = ready_o_1_6[3];
    data_i_1_5[1] = data_o_0_5[2];
    valid_i_1_5[1] = valid_o_0_5[2];
    ready_i_1_5[1] = ready_o_0_5[2];
    data_i_1_5[2] = data_o_2_5[1];
    valid_i_1_5[2] = valid_o_2_5[1];
    ready_i_1_5[2] = ready_o_2_5[1];
    data_i_1_5[0] = data_i[1][5];
    valid_i_1_5[0] = valid_i[1][5];
    ready_i_1_5[0] = ready_i[1][5];
end


/*Router 1,6*/    
merge_router #(
    .input_mask                     (input_mask_1_6),
    .output_sel                     (output_sel_1_6)
)router61(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_1_6),
    .valid_i                        (valid_i_1_6),
    .ready_o                        (ready_o_1_6),
    .data_o                         (data_o_1_6),
    .valid_o                        (valid_o_1_6),
    .ready_i                        (ready_i_1_6)
);


always@(*) begin
    data_i_1_6[3] = data_o_1_5[4];
    valid_i_1_6[3] = valid_o_1_5[4];
    ready_i_1_6[3] = ready_o_1_5[4];
    data_i_1_6[4] = data_o_1_7[3];
    valid_i_1_6[4] = valid_o_1_7[3];
    ready_i_1_6[4] = ready_o_1_7[3];
    data_i_1_6[1] = data_o_0_6[2];
    valid_i_1_6[1] = valid_o_0_6[2];
    ready_i_1_6[1] = ready_o_0_6[2];
    data_i_1_6[2] = data_o_2_6[1];
    valid_i_1_6[2] = valid_o_2_6[1];
    ready_i_1_6[2] = ready_o_2_6[1];
    data_i_1_6[0] = data_i[1][6];
    valid_i_1_6[0] = valid_i[1][6];
    ready_i_1_6[0] = ready_i[1][6];
end


/*Router 1,7*/    
merge_router #(
    .input_mask                     (input_mask_1_7),
    .output_sel                     (output_sel_1_7)
)router71(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_1_7),
    .valid_i                        (valid_i_1_7),
    .ready_o                        (ready_o_1_7),
    .data_o                         (data_o_1_7),
    .valid_o                        (valid_o_1_7),
    .ready_i                        (ready_i_1_7)
);


always@(*) begin
    data_i_1_7[3] = data_o_1_6[4];
    valid_i_1_7[3] = valid_o_1_6[4];
    ready_i_1_7[3] = ready_o_1_6[4];
    data_i_1_7[4] = data_o_1_8[3];
    valid_i_1_7[4] = valid_o_1_8[3];
    ready_i_1_7[4] = ready_o_1_8[3];
    data_i_1_7[1] = data_o_0_7[2];
    valid_i_1_7[1] = valid_o_0_7[2];
    ready_i_1_7[1] = ready_o_0_7[2];
    data_i_1_7[2] = data_o_2_7[1];
    valid_i_1_7[2] = valid_o_2_7[1];
    ready_i_1_7[2] = ready_o_2_7[1];
    data_i_1_7[0] = data_i[1][7];
    valid_i_1_7[0] = valid_i[1][7];
    ready_i_1_7[0] = ready_i[1][7];
end


/*Router 1,8*/    
merge_router #(
    .input_mask                     (input_mask_1_8),
    .output_sel                     (output_sel_1_8)
)router81(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_1_8),
    .valid_i                        (valid_i_1_8),
    .ready_o                        (ready_o_1_8),
    .data_o                         (data_o_1_8),
    .valid_o                        (valid_o_1_8),
    .ready_i                        (ready_i_1_8)
);


always@(*) begin
    data_i_1_8[3] = data_o_1_7[4];
    valid_i_1_8[3] = valid_o_1_7[4];
    ready_i_1_8[3] = ready_o_1_7[4];
    data_i_1_8[4] = data_o_1_9[3];
    valid_i_1_8[4] = valid_o_1_9[3];
    ready_i_1_8[4] = ready_o_1_9[3];
    data_i_1_8[1] = data_o_0_8[2];
    valid_i_1_8[1] = valid_o_0_8[2];
    ready_i_1_8[1] = ready_o_0_8[2];
    data_i_1_8[2] = data_o_2_8[1];
    valid_i_1_8[2] = valid_o_2_8[1];
    ready_i_1_8[2] = ready_o_2_8[1];
    data_i_1_8[0] = data_i[1][8];
    valid_i_1_8[0] = valid_i[1][8];
    ready_i_1_8[0] = ready_i[1][8];
end


/*Router 1,9*/    
merge_router #(
    .input_mask                     (input_mask_1_9),
    .output_sel                     (output_sel_1_9)
)router91(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_1_9),
    .valid_i                        (valid_i_1_9),
    .ready_o                        (ready_o_1_9),
    .data_o                         (data_o_1_9),
    .valid_o                        (valid_o_1_9),
    .ready_i                        (ready_i_1_9)
);


always@(*) begin
    data_i_1_9[3] = data_o_1_8[4];
    valid_i_1_9[3] = valid_o_1_8[4];
    ready_i_1_9[3] = ready_o_1_8[4];
    data_i_1_9[4] = data_o_1_10[3];
    valid_i_1_9[4] = valid_o_1_10[3];
    ready_i_1_9[4] = ready_o_1_10[3];
    data_i_1_9[1] = data_o_0_9[2];
    valid_i_1_9[1] = valid_o_0_9[2];
    ready_i_1_9[1] = ready_o_0_9[2];
    data_i_1_9[2] = data_o_2_9[1];
    valid_i_1_9[2] = valid_o_2_9[1];
    ready_i_1_9[2] = ready_o_2_9[1];
    data_i_1_9[0] = data_i[1][9];
    valid_i_1_9[0] = valid_i[1][9];
    ready_i_1_9[0] = ready_i[1][9];
end


/*Router 1,10*/    
merge_router #(
    .input_mask                     (input_mask_1_10),
    .output_sel                     (output_sel_1_10)
)router101(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_1_10),
    .valid_i                        (valid_i_1_10),
    .ready_o                        (ready_o_1_10),
    .data_o                         (data_o_1_10),
    .valid_o                        (valid_o_1_10),
    .ready_i                        (ready_i_1_10)
);


always@(*) begin
    data_i_1_10[3] = data_o_1_9[4];
    valid_i_1_10[3] = valid_o_1_9[4];
    ready_i_1_10[3] = ready_o_1_9[4];
    data_i_1_10[4] = data_o_1_11[3];
    valid_i_1_10[4] = valid_o_1_11[3];
    ready_i_1_10[4] = ready_o_1_11[3];
    data_i_1_10[1] = data_o_0_10[2];
    valid_i_1_10[1] = valid_o_0_10[2];
    ready_i_1_10[1] = ready_o_0_10[2];
    data_i_1_10[2] = data_o_2_10[1];
    valid_i_1_10[2] = valid_o_2_10[1];
    ready_i_1_10[2] = ready_o_2_10[1];
    data_i_1_10[0] = data_i[1][10];
    valid_i_1_10[0] = valid_i[1][10];
    ready_i_1_10[0] = ready_i[1][10];
end


/*Router 1,11*/    
merge_router #(
    .input_mask                     (input_mask_1_11),
    .output_sel                     (output_sel_1_11)
)router111(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_1_11),
    .valid_i                        (valid_i_1_11),
    .ready_o                        (ready_o_1_11),
    .data_o                         (data_o_1_11),
    .valid_o                        (valid_o_1_11),
    .ready_i                        (ready_i_1_11)
);


always@(*) begin
    data_i_1_11[3] = data_o_1_10[4];
    valid_i_1_11[3] = valid_o_1_10[4];
    ready_i_1_11[3] = ready_o_1_10[4];
    data_i_1_11[4] = data_o_1_12[3];
    valid_i_1_11[4] = valid_o_1_12[3];
    ready_i_1_11[4] = ready_o_1_12[3];
    data_i_1_11[1] = data_o_0_11[2];
    valid_i_1_11[1] = valid_o_0_11[2];
    ready_i_1_11[1] = ready_o_0_11[2];
    data_i_1_11[2] = data_o_2_11[1];
    valid_i_1_11[2] = valid_o_2_11[1];
    ready_i_1_11[2] = ready_o_2_11[1];
    data_i_1_11[0] = data_i[1][11];
    valid_i_1_11[0] = valid_i[1][11];
    ready_i_1_11[0] = ready_i[1][11];
end


/*Router 1,12*/    
merge_router #(
    .input_mask                     (input_mask_1_12),
    .output_sel                     (output_sel_1_12)
)router121(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_1_12),
    .valid_i                        (valid_i_1_12),
    .ready_o                        (ready_o_1_12),
    .data_o                         (data_o_1_12),
    .valid_o                        (valid_o_1_12),
    .ready_i                        (ready_i_1_12)
);


always@(*) begin
    data_i_1_12[3] = data_o_1_11[4];
    valid_i_1_12[3] = valid_o_1_11[4];
    ready_i_1_12[3] = ready_o_1_11[4];
    data_i_1_12[4] = data_o_1_13[3];
    valid_i_1_12[4] = valid_o_1_13[3];
    ready_i_1_12[4] = ready_o_1_13[3];
    data_i_1_12[1] = data_o_0_12[2];
    valid_i_1_12[1] = valid_o_0_12[2];
    ready_i_1_12[1] = ready_o_0_12[2];
    data_i_1_12[2] = data_o_2_12[1];
    valid_i_1_12[2] = valid_o_2_12[1];
    ready_i_1_12[2] = ready_o_2_12[1];
    data_i_1_12[0] = data_i[1][12];
    valid_i_1_12[0] = valid_i[1][12];
    ready_i_1_12[0] = ready_i[1][12];
end


/*Router 1,13*/    
merge_router #(
    .input_mask                     (input_mask_1_13),
    .output_sel                     (output_sel_1_13)
)router131(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_1_13),
    .valid_i                        (valid_i_1_13),
    .ready_o                        (ready_o_1_13),
    .data_o                         (data_o_1_13),
    .valid_o                        (valid_o_1_13),
    .ready_i                        (ready_i_1_13)
);


always@(*) begin
    data_i_1_13[3] = data_o_1_12[4];
    valid_i_1_13[3] = valid_o_1_12[4];
    ready_i_1_13[3] = ready_o_1_12[4];
    data_i_1_13[4] = data_o_1_14[3];
    valid_i_1_13[4] = valid_o_1_14[3];
    ready_i_1_13[4] = ready_o_1_14[3];
    data_i_1_13[1] = data_o_0_13[2];
    valid_i_1_13[1] = valid_o_0_13[2];
    ready_i_1_13[1] = ready_o_0_13[2];
    data_i_1_13[2] = data_o_2_13[1];
    valid_i_1_13[2] = valid_o_2_13[1];
    ready_i_1_13[2] = ready_o_2_13[1];
    data_i_1_13[0] = data_i[1][13];
    valid_i_1_13[0] = valid_i[1][13];
    ready_i_1_13[0] = ready_i[1][13];
end


/*Router 1,14*/    
merge_router #(
    .input_mask                     (input_mask_1_14),
    .output_sel                     (output_sel_1_14)
)router141(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_1_14),
    .valid_i                        (valid_i_1_14),
    .ready_o                        (ready_o_1_14),
    .data_o                         (data_o_1_14),
    .valid_o                        (valid_o_1_14),
    .ready_i                        (ready_i_1_14)
);


always@(*) begin
    data_i_1_14[3] = data_o_1_13[4];
    valid_i_1_14[3] = valid_o_1_13[4];
    ready_i_1_14[3] = ready_o_1_13[4];
    data_i_1_14[4] = data_o_1_15[3];
    valid_i_1_14[4] = valid_o_1_15[3];
    ready_i_1_14[4] = ready_o_1_15[3];
    data_i_1_14[1] = data_o_0_14[2];
    valid_i_1_14[1] = valid_o_0_14[2];
    ready_i_1_14[1] = ready_o_0_14[2];
    data_i_1_14[2] = data_o_2_14[1];
    valid_i_1_14[2] = valid_o_2_14[1];
    ready_i_1_14[2] = ready_o_2_14[1];
    data_i_1_14[0] = data_i[1][14];
    valid_i_1_14[0] = valid_i[1][14];
    ready_i_1_14[0] = ready_i[1][14];
end


/*Router 1,15*/    
merge_router #(
    .input_mask                     (input_mask_1_15),
    .output_sel                     (output_sel_1_15)
)router151(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_1_15),
    .valid_i                        (valid_i_1_15),
    .ready_o                        (ready_o_1_15),
    .data_o                         (data_o_1_15),
    .valid_o                        (valid_o_1_15),
    .ready_i                        (ready_i_1_15)
);


always@(*) begin
    data_i_1_15[3] = data_o_1_14[4];
    valid_i_1_15[3] = valid_o_1_14[4];
    ready_i_1_15[3] = ready_o_1_14[4];
    data_i_1_15[4] = data_o_1_16[3];
    valid_i_1_15[4] = valid_o_1_16[3];
    ready_i_1_15[4] = ready_o_1_16[3];
    data_i_1_15[1] = data_o_0_15[2];
    valid_i_1_15[1] = valid_o_0_15[2];
    ready_i_1_15[1] = ready_o_0_15[2];
    data_i_1_15[2] = data_o_2_15[1];
    valid_i_1_15[2] = valid_o_2_15[1];
    ready_i_1_15[2] = ready_o_2_15[1];
    data_i_1_15[0] = data_i[1][15];
    valid_i_1_15[0] = valid_i[1][15];
    ready_i_1_15[0] = ready_i[1][15];
end


/*Router 1,16*/    
merge_router #(
    .input_mask                     (input_mask_1_16),
    .output_sel                     (output_sel_1_16)
)router161(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_1_16),
    .valid_i                        (valid_i_1_16),
    .ready_o                        (ready_o_1_16),
    .data_o                         (data_o_1_16),
    .valid_o                        (valid_o_1_16),
    .ready_i                        (ready_i_1_16)
);


always@(*) begin
    data_i_1_16[3] = data_o_1_15[4];
    valid_i_1_16[3] = valid_o_1_15[4];
    ready_i_1_16[3] = ready_o_1_15[4];
    data_i_1_16[4] = data_o_1_17[3];
    valid_i_1_16[4] = valid_o_1_17[3];
    ready_i_1_16[4] = ready_o_1_17[3];
    data_i_1_16[1] = data_o_0_16[2];
    valid_i_1_16[1] = valid_o_0_16[2];
    ready_i_1_16[1] = ready_o_0_16[2];
    data_i_1_16[2] = data_o_2_16[1];
    valid_i_1_16[2] = valid_o_2_16[1];
    ready_i_1_16[2] = ready_o_2_16[1];
    data_i_1_16[0] = data_i[1][16];
    valid_i_1_16[0] = valid_i[1][16];
    ready_i_1_16[0] = ready_i[1][16];
end


/*Router 1,17*/    
merge_router #(
    .input_mask                     (input_mask_1_17),
    .output_sel                     (output_sel_1_17)
)router171(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_1_17),
    .valid_i                        (valid_i_1_17),
    .ready_o                        (ready_o_1_17),
    .data_o                         (data_o_1_17),
    .valid_o                        (valid_o_1_17),
    .ready_i                        (ready_i_1_17)
);


always@(*) begin
    data_i_1_17[3] = data_o_1_16[4];
    valid_i_1_17[3] = valid_o_1_16[4];
    ready_i_1_17[3] = ready_o_1_16[4];
    data_i_1_17[4] = data_o_1_18[3];
    valid_i_1_17[4] = valid_o_1_18[3];
    ready_i_1_17[4] = ready_o_1_18[3];
    data_i_1_17[1] = data_o_0_17[2];
    valid_i_1_17[1] = valid_o_0_17[2];
    ready_i_1_17[1] = ready_o_0_17[2];
    data_i_1_17[2] = data_o_2_17[1];
    valid_i_1_17[2] = valid_o_2_17[1];
    ready_i_1_17[2] = ready_o_2_17[1];
    data_i_1_17[0] = data_i[1][17];
    valid_i_1_17[0] = valid_i[1][17];
    ready_i_1_17[0] = ready_i[1][17];
end


/*Router 1,18*/    
merge_router #(
    .input_mask                     (input_mask_1_18),
    .output_sel                     (output_sel_1_18)
)router181(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_1_18),
    .valid_i                        (valid_i_1_18),
    .ready_o                        (ready_o_1_18),
    .data_o                         (data_o_1_18),
    .valid_o                        (valid_o_1_18),
    .ready_i                        (ready_i_1_18)
);


always@(*) begin
    data_i_1_18[3] = data_o_1_17[4];
    valid_i_1_18[3] = valid_o_1_17[4];
    ready_i_1_18[3] = ready_o_1_17[4];
    data_i_1_18[4] = data_o_1_19[3];
    valid_i_1_18[4] = valid_o_1_19[3];
    ready_i_1_18[4] = ready_o_1_19[3];
    data_i_1_18[1] = data_o_0_18[2];
    valid_i_1_18[1] = valid_o_0_18[2];
    ready_i_1_18[1] = ready_o_0_18[2];
    data_i_1_18[2] = data_o_2_18[1];
    valid_i_1_18[2] = valid_o_2_18[1];
    ready_i_1_18[2] = ready_o_2_18[1];
    data_i_1_18[0] = data_i[1][18];
    valid_i_1_18[0] = valid_i[1][18];
    ready_i_1_18[0] = ready_i[1][18];
end


/*Router 1,19*/    
merge_router #(
    .input_mask                     (input_mask_1_19),
    .output_sel                     (output_sel_1_19)
)router191(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_1_19),
    .valid_i                        (valid_i_1_19),
    .ready_o                        (ready_o_1_19),
    .data_o                         (data_o_1_19),
    .valid_o                        (valid_o_1_19),
    .ready_i                        (ready_i_1_19)
);


always@(*) begin
    data_i_1_19[3] = data_o_1_18[4];
    valid_i_1_19[3] = valid_o_1_18[4];
    ready_i_1_19[3] = ready_o_1_18[4];
    data_i_1_19[4] = data_o_1_20[3];
    valid_i_1_19[4] = valid_o_1_20[3];
    ready_i_1_19[4] = ready_o_1_20[3];
    data_i_1_19[1] = data_o_0_19[2];
    valid_i_1_19[1] = valid_o_0_19[2];
    ready_i_1_19[1] = ready_o_0_19[2];
    data_i_1_19[2] = data_o_2_19[1];
    valid_i_1_19[2] = valid_o_2_19[1];
    ready_i_1_19[2] = ready_o_2_19[1];
    data_i_1_19[0] = data_i[1][19];
    valid_i_1_19[0] = valid_i[1][19];
    ready_i_1_19[0] = ready_i[1][19];
end


/*Router 1,20*/    
merge_router #(
    .input_mask                     (input_mask_1_20),
    .output_sel                     (output_sel_1_20)
)router201(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_1_20),
    .valid_i                        (valid_i_1_20),
    .ready_o                        (ready_o_1_20),
    .data_o                         (data_o_1_20),
    .valid_o                        (valid_o_1_20),
    .ready_i                        (ready_i_1_20)
);


always@(*) begin
    data_i_1_20[3] = data_o_1_19[4];
    valid_i_1_20[3] = valid_o_1_19[4];
    ready_i_1_20[3] = ready_o_1_19[4];
    data_i_1_20[4] = data_o_1_21[3];
    valid_i_1_20[4] = valid_o_1_21[3];
    ready_i_1_20[4] = ready_o_1_21[3];
    data_i_1_20[1] = data_o_0_20[2];
    valid_i_1_20[1] = valid_o_0_20[2];
    ready_i_1_20[1] = ready_o_0_20[2];
    data_i_1_20[2] = data_o_2_20[1];
    valid_i_1_20[2] = valid_o_2_20[1];
    ready_i_1_20[2] = ready_o_2_20[1];
    data_i_1_20[0] = data_i[1][20];
    valid_i_1_20[0] = valid_i[1][20];
    ready_i_1_20[0] = ready_i[1][20];
end


/*Router 1,21*/    
merge_router #(
    .input_mask                     (input_mask_1_21),
    .output_sel                     (output_sel_1_21)
)router211(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_1_21),
    .valid_i                        (valid_i_1_21),
    .ready_o                        (ready_o_1_21),
    .data_o                         (data_o_1_21),
    .valid_o                        (valid_o_1_21),
    .ready_i                        (ready_i_1_21)
);


always@(*) begin
    data_i_1_21[3] = data_o_1_20[4];
    valid_i_1_21[3] = valid_o_1_20[4];
    ready_i_1_21[3] = ready_o_1_20[4];
    data_i_1_21[4] = data_o_1_22[3];
    valid_i_1_21[4] = valid_o_1_22[3];
    ready_i_1_21[4] = ready_o_1_22[3];
    data_i_1_21[1] = data_o_0_21[2];
    valid_i_1_21[1] = valid_o_0_21[2];
    ready_i_1_21[1] = ready_o_0_21[2];
    data_i_1_21[2] = data_o_2_21[1];
    valid_i_1_21[2] = valid_o_2_21[1];
    ready_i_1_21[2] = ready_o_2_21[1];
    data_i_1_21[0] = data_i[1][21];
    valid_i_1_21[0] = valid_i[1][21];
    ready_i_1_21[0] = ready_i[1][21];
end


/*Router 1,22*/    
merge_router #(
    .input_mask                     (input_mask_1_22),
    .output_sel                     (output_sel_1_22)
)router221(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_1_22),
    .valid_i                        (valid_i_1_22),
    .ready_o                        (ready_o_1_22),
    .data_o                         (data_o_1_22),
    .valid_o                        (valid_o_1_22),
    .ready_i                        (ready_i_1_22)
);


always@(*) begin
    data_i_1_22[3] = data_o_1_21[4];
    valid_i_1_22[3] = valid_o_1_21[4];
    ready_i_1_22[3] = ready_o_1_21[4];
    data_i_1_22[4] = data_o_1_23[3];
    valid_i_1_22[4] = valid_o_1_23[3];
    ready_i_1_22[4] = ready_o_1_23[3];
    data_i_1_22[1] = data_o_0_22[2];
    valid_i_1_22[1] = valid_o_0_22[2];
    ready_i_1_22[1] = ready_o_0_22[2];
    data_i_1_22[2] = data_o_2_22[1];
    valid_i_1_22[2] = valid_o_2_22[1];
    ready_i_1_22[2] = ready_o_2_22[1];
    data_i_1_22[0] = data_i[1][22];
    valid_i_1_22[0] = valid_i[1][22];
    ready_i_1_22[0] = ready_i[1][22];
end


/*Router 1,23*/    
merge_router #(
    .input_mask                     (input_mask_1_23),
    .output_sel                     (output_sel_1_23)
)router231(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_1_23),
    .valid_i                        (valid_i_1_23),
    .ready_o                        (ready_o_1_23),
    .data_o                         (data_o_1_23),
    .valid_o                        (valid_o_1_23),
    .ready_i                        (ready_i_1_23)
);


always@(*) begin
    data_i_1_23[3] = data_o_1_22[4];
    valid_i_1_23[3] = valid_o_1_22[4];
    ready_i_1_23[3] = ready_o_1_22[4];
    data_i_1_23[4] = data_o_1_24[3];
    valid_i_1_23[4] = valid_o_1_24[3];
    ready_i_1_23[4] = ready_o_1_24[3];
    data_i_1_23[1] = data_o_0_23[2];
    valid_i_1_23[1] = valid_o_0_23[2];
    ready_i_1_23[1] = ready_o_0_23[2];
    data_i_1_23[2] = data_o_2_23[1];
    valid_i_1_23[2] = valid_o_2_23[1];
    ready_i_1_23[2] = ready_o_2_23[1];
    data_i_1_23[0] = data_i[1][23];
    valid_i_1_23[0] = valid_i[1][23];
    ready_i_1_23[0] = ready_i[1][23];
end


/*Router 1,24*/    
merge_router #(
    .input_mask                     (input_mask_1_24),
    .output_sel                     (output_sel_1_24)
)router241(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_1_24),
    .valid_i                        (valid_i_1_24),
    .ready_o                        (ready_o_1_24),
    .data_o                         (data_o_1_24),
    .valid_o                        (valid_o_1_24),
    .ready_i                        (ready_i_1_24)
);


always@(*) begin
    data_i_1_24[3] = data_o_1_23[4];
    valid_i_1_24[3] = valid_o_1_23[4];
    ready_i_1_24[3] = ready_o_1_23[4];
    data_i_1_24[1] = data_o_0_24[2];
    valid_i_1_24[1] = valid_o_0_24[2];
    ready_i_1_24[1] = ready_o_0_24[2];
    data_i_1_24[2] = data_o_2_24[1];
    valid_i_1_24[2] = valid_o_2_24[1];
    ready_i_1_24[2] = ready_o_2_24[1];
    data_i_1_24[0] = data_i[1][24];
    valid_i_1_24[0] = valid_i[1][24];
    ready_i_1_24[0] = ready_i[1][24];
end


/*Router 2,0*/    
merge_router #(
    .input_mask                     (input_mask_2_0),
    .output_sel                     (output_sel_2_0)
)router2(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_2_0),
    .valid_i                        (valid_i_2_0),
    .ready_o                        (ready_o_2_0),
    .data_o                         (data_o_2_0),
    .valid_o                        (valid_o_2_0),
    .ready_i                        (ready_i_2_0)
);


always@(*) begin
    data_i_2_0[4] = data_o_2_1[3];
    valid_i_2_0[4] = valid_o_2_1[3];
    ready_i_2_0[4] = ready_o_2_1[3];
    data_i_2_0[1] = data_o_1_0[2];
    valid_i_2_0[1] = valid_o_1_0[2];
    ready_i_2_0[1] = ready_o_1_0[2];
    data_i_2_0[2] = data_o_3_0[1];
    valid_i_2_0[2] = valid_o_3_0[1];
    ready_i_2_0[2] = ready_o_3_0[1];
    data_i_2_0[0] = data_i[2][0];
    valid_i_2_0[0] = valid_i[2][0];
    ready_i_2_0[0] = ready_i[2][0];
end


/*Router 2,1*/    
merge_router #(
    .input_mask                     (input_mask_2_1),
    .output_sel                     (output_sel_2_1)
)router12(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_2_1),
    .valid_i                        (valid_i_2_1),
    .ready_o                        (ready_o_2_1),
    .data_o                         (data_o_2_1),
    .valid_o                        (valid_o_2_1),
    .ready_i                        (ready_i_2_1)
);


always@(*) begin
    data_i_2_1[3] = data_o_2_0[4];
    valid_i_2_1[3] = valid_o_2_0[4];
    ready_i_2_1[3] = ready_o_2_0[4];
    data_i_2_1[4] = data_o_2_2[3];
    valid_i_2_1[4] = valid_o_2_2[3];
    ready_i_2_1[4] = ready_o_2_2[3];
    data_i_2_1[1] = data_o_1_1[2];
    valid_i_2_1[1] = valid_o_1_1[2];
    ready_i_2_1[1] = ready_o_1_1[2];
    data_i_2_1[2] = data_o_3_1[1];
    valid_i_2_1[2] = valid_o_3_1[1];
    ready_i_2_1[2] = ready_o_3_1[1];
    data_i_2_1[0] = data_i[2][1];
    valid_i_2_1[0] = valid_i[2][1];
    ready_i_2_1[0] = ready_i[2][1];
end


/*Router 2,2*/    
merge_router #(
    .input_mask                     (input_mask_2_2),
    .output_sel                     (output_sel_2_2)
)router22(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_2_2),
    .valid_i                        (valid_i_2_2),
    .ready_o                        (ready_o_2_2),
    .data_o                         (data_o_2_2),
    .valid_o                        (valid_o_2_2),
    .ready_i                        (ready_i_2_2)
);


always@(*) begin
    data_i_2_2[3] = data_o_2_1[4];
    valid_i_2_2[3] = valid_o_2_1[4];
    ready_i_2_2[3] = ready_o_2_1[4];
    data_i_2_2[4] = data_o_2_3[3];
    valid_i_2_2[4] = valid_o_2_3[3];
    ready_i_2_2[4] = ready_o_2_3[3];
    data_i_2_2[1] = data_o_1_2[2];
    valid_i_2_2[1] = valid_o_1_2[2];
    ready_i_2_2[1] = ready_o_1_2[2];
    data_i_2_2[2] = data_o_3_2[1];
    valid_i_2_2[2] = valid_o_3_2[1];
    ready_i_2_2[2] = ready_o_3_2[1];
    data_i_2_2[0] = data_i[2][2];
    valid_i_2_2[0] = valid_i[2][2];
    ready_i_2_2[0] = ready_i[2][2];
end


/*Router 2,3*/    
merge_router #(
    .input_mask                     (input_mask_2_3),
    .output_sel                     (output_sel_2_3)
)router32(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_2_3),
    .valid_i                        (valid_i_2_3),
    .ready_o                        (ready_o_2_3),
    .data_o                         (data_o_2_3),
    .valid_o                        (valid_o_2_3),
    .ready_i                        (ready_i_2_3)
);


always@(*) begin
    data_i_2_3[3] = data_o_2_2[4];
    valid_i_2_3[3] = valid_o_2_2[4];
    ready_i_2_3[3] = ready_o_2_2[4];
    data_i_2_3[4] = data_o_2_4[3];
    valid_i_2_3[4] = valid_o_2_4[3];
    ready_i_2_3[4] = ready_o_2_4[3];
    data_i_2_3[1] = data_o_1_3[2];
    valid_i_2_3[1] = valid_o_1_3[2];
    ready_i_2_3[1] = ready_o_1_3[2];
    data_i_2_3[2] = data_o_3_3[1];
    valid_i_2_3[2] = valid_o_3_3[1];
    ready_i_2_3[2] = ready_o_3_3[1];
    data_i_2_3[0] = data_i[2][3];
    valid_i_2_3[0] = valid_i[2][3];
    ready_i_2_3[0] = ready_i[2][3];
end


/*Router 2,4*/    
merge_router #(
    .input_mask                     (input_mask_2_4),
    .output_sel                     (output_sel_2_4)
)router42(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_2_4),
    .valid_i                        (valid_i_2_4),
    .ready_o                        (ready_o_2_4),
    .data_o                         (data_o_2_4),
    .valid_o                        (valid_o_2_4),
    .ready_i                        (ready_i_2_4)
);


always@(*) begin
    data_i_2_4[3] = data_o_2_3[4];
    valid_i_2_4[3] = valid_o_2_3[4];
    ready_i_2_4[3] = ready_o_2_3[4];
    data_i_2_4[4] = data_o_2_5[3];
    valid_i_2_4[4] = valid_o_2_5[3];
    ready_i_2_4[4] = ready_o_2_5[3];
    data_i_2_4[1] = data_o_1_4[2];
    valid_i_2_4[1] = valid_o_1_4[2];
    ready_i_2_4[1] = ready_o_1_4[2];
    data_i_2_4[2] = data_o_3_4[1];
    valid_i_2_4[2] = valid_o_3_4[1];
    ready_i_2_4[2] = ready_o_3_4[1];
    data_i_2_4[0] = data_i[2][4];
    valid_i_2_4[0] = valid_i[2][4];
    ready_i_2_4[0] = ready_i[2][4];
end


/*Router 2,5*/    
merge_router #(
    .input_mask                     (input_mask_2_5),
    .output_sel                     (output_sel_2_5)
)router52(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_2_5),
    .valid_i                        (valid_i_2_5),
    .ready_o                        (ready_o_2_5),
    .data_o                         (data_o_2_5),
    .valid_o                        (valid_o_2_5),
    .ready_i                        (ready_i_2_5)
);


always@(*) begin
    data_i_2_5[3] = data_o_2_4[4];
    valid_i_2_5[3] = valid_o_2_4[4];
    ready_i_2_5[3] = ready_o_2_4[4];
    data_i_2_5[4] = data_o_2_6[3];
    valid_i_2_5[4] = valid_o_2_6[3];
    ready_i_2_5[4] = ready_o_2_6[3];
    data_i_2_5[1] = data_o_1_5[2];
    valid_i_2_5[1] = valid_o_1_5[2];
    ready_i_2_5[1] = ready_o_1_5[2];
    data_i_2_5[2] = data_o_3_5[1];
    valid_i_2_5[2] = valid_o_3_5[1];
    ready_i_2_5[2] = ready_o_3_5[1];
    data_i_2_5[0] = data_i[2][5];
    valid_i_2_5[0] = valid_i[2][5];
    ready_i_2_5[0] = ready_i[2][5];
end


/*Router 2,6*/    
merge_router #(
    .input_mask                     (input_mask_2_6),
    .output_sel                     (output_sel_2_6)
)router62(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_2_6),
    .valid_i                        (valid_i_2_6),
    .ready_o                        (ready_o_2_6),
    .data_o                         (data_o_2_6),
    .valid_o                        (valid_o_2_6),
    .ready_i                        (ready_i_2_6)
);


always@(*) begin
    data_i_2_6[3] = data_o_2_5[4];
    valid_i_2_6[3] = valid_o_2_5[4];
    ready_i_2_6[3] = ready_o_2_5[4];
    data_i_2_6[4] = data_o_2_7[3];
    valid_i_2_6[4] = valid_o_2_7[3];
    ready_i_2_6[4] = ready_o_2_7[3];
    data_i_2_6[1] = data_o_1_6[2];
    valid_i_2_6[1] = valid_o_1_6[2];
    ready_i_2_6[1] = ready_o_1_6[2];
    data_i_2_6[2] = data_o_3_6[1];
    valid_i_2_6[2] = valid_o_3_6[1];
    ready_i_2_6[2] = ready_o_3_6[1];
    data_i_2_6[0] = data_i[2][6];
    valid_i_2_6[0] = valid_i[2][6];
    ready_i_2_6[0] = ready_i[2][6];
end


/*Router 2,7*/    
merge_router #(
    .input_mask                     (input_mask_2_7),
    .output_sel                     (output_sel_2_7)
)router72(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_2_7),
    .valid_i                        (valid_i_2_7),
    .ready_o                        (ready_o_2_7),
    .data_o                         (data_o_2_7),
    .valid_o                        (valid_o_2_7),
    .ready_i                        (ready_i_2_7)
);


always@(*) begin
    data_i_2_7[3] = data_o_2_6[4];
    valid_i_2_7[3] = valid_o_2_6[4];
    ready_i_2_7[3] = ready_o_2_6[4];
    data_i_2_7[4] = data_o_2_8[3];
    valid_i_2_7[4] = valid_o_2_8[3];
    ready_i_2_7[4] = ready_o_2_8[3];
    data_i_2_7[1] = data_o_1_7[2];
    valid_i_2_7[1] = valid_o_1_7[2];
    ready_i_2_7[1] = ready_o_1_7[2];
    data_i_2_7[2] = data_o_3_7[1];
    valid_i_2_7[2] = valid_o_3_7[1];
    ready_i_2_7[2] = ready_o_3_7[1];
    data_i_2_7[0] = data_i[2][7];
    valid_i_2_7[0] = valid_i[2][7];
    ready_i_2_7[0] = ready_i[2][7];
end


/*Router 2,8*/    
merge_router #(
    .input_mask                     (input_mask_2_8),
    .output_sel                     (output_sel_2_8)
)router82(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_2_8),
    .valid_i                        (valid_i_2_8),
    .ready_o                        (ready_o_2_8),
    .data_o                         (data_o_2_8),
    .valid_o                        (valid_o_2_8),
    .ready_i                        (ready_i_2_8)
);


always@(*) begin
    data_i_2_8[3] = data_o_2_7[4];
    valid_i_2_8[3] = valid_o_2_7[4];
    ready_i_2_8[3] = ready_o_2_7[4];
    data_i_2_8[4] = data_o_2_9[3];
    valid_i_2_8[4] = valid_o_2_9[3];
    ready_i_2_8[4] = ready_o_2_9[3];
    data_i_2_8[1] = data_o_1_8[2];
    valid_i_2_8[1] = valid_o_1_8[2];
    ready_i_2_8[1] = ready_o_1_8[2];
    data_i_2_8[2] = data_o_3_8[1];
    valid_i_2_8[2] = valid_o_3_8[1];
    ready_i_2_8[2] = ready_o_3_8[1];
    data_i_2_8[0] = data_i[2][8];
    valid_i_2_8[0] = valid_i[2][8];
    ready_i_2_8[0] = ready_i[2][8];
end


/*Router 2,9*/    
merge_router #(
    .input_mask                     (input_mask_2_9),
    .output_sel                     (output_sel_2_9)
)router92(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_2_9),
    .valid_i                        (valid_i_2_9),
    .ready_o                        (ready_o_2_9),
    .data_o                         (data_o_2_9),
    .valid_o                        (valid_o_2_9),
    .ready_i                        (ready_i_2_9)
);


always@(*) begin
    data_i_2_9[3] = data_o_2_8[4];
    valid_i_2_9[3] = valid_o_2_8[4];
    ready_i_2_9[3] = ready_o_2_8[4];
    data_i_2_9[4] = data_o_2_10[3];
    valid_i_2_9[4] = valid_o_2_10[3];
    ready_i_2_9[4] = ready_o_2_10[3];
    data_i_2_9[1] = data_o_1_9[2];
    valid_i_2_9[1] = valid_o_1_9[2];
    ready_i_2_9[1] = ready_o_1_9[2];
    data_i_2_9[2] = data_o_3_9[1];
    valid_i_2_9[2] = valid_o_3_9[1];
    ready_i_2_9[2] = ready_o_3_9[1];
    data_i_2_9[0] = data_i[2][9];
    valid_i_2_9[0] = valid_i[2][9];
    ready_i_2_9[0] = ready_i[2][9];
end


/*Router 2,10*/    
merge_router #(
    .input_mask                     (input_mask_2_10),
    .output_sel                     (output_sel_2_10)
)router102(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_2_10),
    .valid_i                        (valid_i_2_10),
    .ready_o                        (ready_o_2_10),
    .data_o                         (data_o_2_10),
    .valid_o                        (valid_o_2_10),
    .ready_i                        (ready_i_2_10)
);


always@(*) begin
    data_i_2_10[3] = data_o_2_9[4];
    valid_i_2_10[3] = valid_o_2_9[4];
    ready_i_2_10[3] = ready_o_2_9[4];
    data_i_2_10[4] = data_o_2_11[3];
    valid_i_2_10[4] = valid_o_2_11[3];
    ready_i_2_10[4] = ready_o_2_11[3];
    data_i_2_10[1] = data_o_1_10[2];
    valid_i_2_10[1] = valid_o_1_10[2];
    ready_i_2_10[1] = ready_o_1_10[2];
    data_i_2_10[2] = data_o_3_10[1];
    valid_i_2_10[2] = valid_o_3_10[1];
    ready_i_2_10[2] = ready_o_3_10[1];
    data_i_2_10[0] = data_i[2][10];
    valid_i_2_10[0] = valid_i[2][10];
    ready_i_2_10[0] = ready_i[2][10];
end


/*Router 2,11*/    
merge_router #(
    .input_mask                     (input_mask_2_11),
    .output_sel                     (output_sel_2_11)
)router112(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_2_11),
    .valid_i                        (valid_i_2_11),
    .ready_o                        (ready_o_2_11),
    .data_o                         (data_o_2_11),
    .valid_o                        (valid_o_2_11),
    .ready_i                        (ready_i_2_11)
);


always@(*) begin
    data_i_2_11[3] = data_o_2_10[4];
    valid_i_2_11[3] = valid_o_2_10[4];
    ready_i_2_11[3] = ready_o_2_10[4];
    data_i_2_11[4] = data_o_2_12[3];
    valid_i_2_11[4] = valid_o_2_12[3];
    ready_i_2_11[4] = ready_o_2_12[3];
    data_i_2_11[1] = data_o_1_11[2];
    valid_i_2_11[1] = valid_o_1_11[2];
    ready_i_2_11[1] = ready_o_1_11[2];
    data_i_2_11[2] = data_o_3_11[1];
    valid_i_2_11[2] = valid_o_3_11[1];
    ready_i_2_11[2] = ready_o_3_11[1];
    data_i_2_11[0] = data_i[2][11];
    valid_i_2_11[0] = valid_i[2][11];
    ready_i_2_11[0] = ready_i[2][11];
end


/*Router 2,12*/    
merge_router #(
    .input_mask                     (input_mask_2_12),
    .output_sel                     (output_sel_2_12)
)router122(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_2_12),
    .valid_i                        (valid_i_2_12),
    .ready_o                        (ready_o_2_12),
    .data_o                         (data_o_2_12),
    .valid_o                        (valid_o_2_12),
    .ready_i                        (ready_i_2_12)
);


always@(*) begin
    data_i_2_12[3] = data_o_2_11[4];
    valid_i_2_12[3] = valid_o_2_11[4];
    ready_i_2_12[3] = ready_o_2_11[4];
    data_i_2_12[4] = data_o_2_13[3];
    valid_i_2_12[4] = valid_o_2_13[3];
    ready_i_2_12[4] = ready_o_2_13[3];
    data_i_2_12[1] = data_o_1_12[2];
    valid_i_2_12[1] = valid_o_1_12[2];
    ready_i_2_12[1] = ready_o_1_12[2];
    data_i_2_12[2] = data_o_3_12[1];
    valid_i_2_12[2] = valid_o_3_12[1];
    ready_i_2_12[2] = ready_o_3_12[1];
    data_i_2_12[0] = data_i[2][12];
    valid_i_2_12[0] = valid_i[2][12];
    ready_i_2_12[0] = ready_i[2][12];
end


/*Router 2,13*/    
merge_router #(
    .input_mask                     (input_mask_2_13),
    .output_sel                     (output_sel_2_13)
)router132(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_2_13),
    .valid_i                        (valid_i_2_13),
    .ready_o                        (ready_o_2_13),
    .data_o                         (data_o_2_13),
    .valid_o                        (valid_o_2_13),
    .ready_i                        (ready_i_2_13)
);


always@(*) begin
    data_i_2_13[3] = data_o_2_12[4];
    valid_i_2_13[3] = valid_o_2_12[4];
    ready_i_2_13[3] = ready_o_2_12[4];
    data_i_2_13[4] = data_o_2_14[3];
    valid_i_2_13[4] = valid_o_2_14[3];
    ready_i_2_13[4] = ready_o_2_14[3];
    data_i_2_13[1] = data_o_1_13[2];
    valid_i_2_13[1] = valid_o_1_13[2];
    ready_i_2_13[1] = ready_o_1_13[2];
    data_i_2_13[2] = data_o_3_13[1];
    valid_i_2_13[2] = valid_o_3_13[1];
    ready_i_2_13[2] = ready_o_3_13[1];
    data_i_2_13[0] = data_i[2][13];
    valid_i_2_13[0] = valid_i[2][13];
    ready_i_2_13[0] = ready_i[2][13];
end


/*Router 2,14*/    
merge_router #(
    .input_mask                     (input_mask_2_14),
    .output_sel                     (output_sel_2_14)
)router142(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_2_14),
    .valid_i                        (valid_i_2_14),
    .ready_o                        (ready_o_2_14),
    .data_o                         (data_o_2_14),
    .valid_o                        (valid_o_2_14),
    .ready_i                        (ready_i_2_14)
);


always@(*) begin
    data_i_2_14[3] = data_o_2_13[4];
    valid_i_2_14[3] = valid_o_2_13[4];
    ready_i_2_14[3] = ready_o_2_13[4];
    data_i_2_14[4] = data_o_2_15[3];
    valid_i_2_14[4] = valid_o_2_15[3];
    ready_i_2_14[4] = ready_o_2_15[3];
    data_i_2_14[1] = data_o_1_14[2];
    valid_i_2_14[1] = valid_o_1_14[2];
    ready_i_2_14[1] = ready_o_1_14[2];
    data_i_2_14[2] = data_o_3_14[1];
    valid_i_2_14[2] = valid_o_3_14[1];
    ready_i_2_14[2] = ready_o_3_14[1];
    data_i_2_14[0] = data_i[2][14];
    valid_i_2_14[0] = valid_i[2][14];
    ready_i_2_14[0] = ready_i[2][14];
end


/*Router 2,15*/    
merge_router #(
    .input_mask                     (input_mask_2_15),
    .output_sel                     (output_sel_2_15)
)router152(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_2_15),
    .valid_i                        (valid_i_2_15),
    .ready_o                        (ready_o_2_15),
    .data_o                         (data_o_2_15),
    .valid_o                        (valid_o_2_15),
    .ready_i                        (ready_i_2_15)
);


always@(*) begin
    data_i_2_15[3] = data_o_2_14[4];
    valid_i_2_15[3] = valid_o_2_14[4];
    ready_i_2_15[3] = ready_o_2_14[4];
    data_i_2_15[4] = data_o_2_16[3];
    valid_i_2_15[4] = valid_o_2_16[3];
    ready_i_2_15[4] = ready_o_2_16[3];
    data_i_2_15[1] = data_o_1_15[2];
    valid_i_2_15[1] = valid_o_1_15[2];
    ready_i_2_15[1] = ready_o_1_15[2];
    data_i_2_15[2] = data_o_3_15[1];
    valid_i_2_15[2] = valid_o_3_15[1];
    ready_i_2_15[2] = ready_o_3_15[1];
    data_i_2_15[0] = data_i[2][15];
    valid_i_2_15[0] = valid_i[2][15];
    ready_i_2_15[0] = ready_i[2][15];
end


/*Router 2,16*/    
merge_router #(
    .input_mask                     (input_mask_2_16),
    .output_sel                     (output_sel_2_16)
)router162(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_2_16),
    .valid_i                        (valid_i_2_16),
    .ready_o                        (ready_o_2_16),
    .data_o                         (data_o_2_16),
    .valid_o                        (valid_o_2_16),
    .ready_i                        (ready_i_2_16)
);


always@(*) begin
    data_i_2_16[3] = data_o_2_15[4];
    valid_i_2_16[3] = valid_o_2_15[4];
    ready_i_2_16[3] = ready_o_2_15[4];
    data_i_2_16[4] = data_o_2_17[3];
    valid_i_2_16[4] = valid_o_2_17[3];
    ready_i_2_16[4] = ready_o_2_17[3];
    data_i_2_16[1] = data_o_1_16[2];
    valid_i_2_16[1] = valid_o_1_16[2];
    ready_i_2_16[1] = ready_o_1_16[2];
    data_i_2_16[2] = data_o_3_16[1];
    valid_i_2_16[2] = valid_o_3_16[1];
    ready_i_2_16[2] = ready_o_3_16[1];
    data_i_2_16[0] = data_i[2][16];
    valid_i_2_16[0] = valid_i[2][16];
    ready_i_2_16[0] = ready_i[2][16];
end


/*Router 2,17*/    
merge_router #(
    .input_mask                     (input_mask_2_17),
    .output_sel                     (output_sel_2_17)
)router172(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_2_17),
    .valid_i                        (valid_i_2_17),
    .ready_o                        (ready_o_2_17),
    .data_o                         (data_o_2_17),
    .valid_o                        (valid_o_2_17),
    .ready_i                        (ready_i_2_17)
);


always@(*) begin
    data_i_2_17[3] = data_o_2_16[4];
    valid_i_2_17[3] = valid_o_2_16[4];
    ready_i_2_17[3] = ready_o_2_16[4];
    data_i_2_17[4] = data_o_2_18[3];
    valid_i_2_17[4] = valid_o_2_18[3];
    ready_i_2_17[4] = ready_o_2_18[3];
    data_i_2_17[1] = data_o_1_17[2];
    valid_i_2_17[1] = valid_o_1_17[2];
    ready_i_2_17[1] = ready_o_1_17[2];
    data_i_2_17[2] = data_o_3_17[1];
    valid_i_2_17[2] = valid_o_3_17[1];
    ready_i_2_17[2] = ready_o_3_17[1];
    data_i_2_17[0] = data_i[2][17];
    valid_i_2_17[0] = valid_i[2][17];
    ready_i_2_17[0] = ready_i[2][17];
end


/*Router 2,18*/    
merge_router #(
    .input_mask                     (input_mask_2_18),
    .output_sel                     (output_sel_2_18)
)router182(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_2_18),
    .valid_i                        (valid_i_2_18),
    .ready_o                        (ready_o_2_18),
    .data_o                         (data_o_2_18),
    .valid_o                        (valid_o_2_18),
    .ready_i                        (ready_i_2_18)
);


always@(*) begin
    data_i_2_18[3] = data_o_2_17[4];
    valid_i_2_18[3] = valid_o_2_17[4];
    ready_i_2_18[3] = ready_o_2_17[4];
    data_i_2_18[4] = data_o_2_19[3];
    valid_i_2_18[4] = valid_o_2_19[3];
    ready_i_2_18[4] = ready_o_2_19[3];
    data_i_2_18[1] = data_o_1_18[2];
    valid_i_2_18[1] = valid_o_1_18[2];
    ready_i_2_18[1] = ready_o_1_18[2];
    data_i_2_18[2] = data_o_3_18[1];
    valid_i_2_18[2] = valid_o_3_18[1];
    ready_i_2_18[2] = ready_o_3_18[1];
    data_i_2_18[0] = data_i[2][18];
    valid_i_2_18[0] = valid_i[2][18];
    ready_i_2_18[0] = ready_i[2][18];
end


/*Router 2,19*/    
merge_router #(
    .input_mask                     (input_mask_2_19),
    .output_sel                     (output_sel_2_19)
)router192(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_2_19),
    .valid_i                        (valid_i_2_19),
    .ready_o                        (ready_o_2_19),
    .data_o                         (data_o_2_19),
    .valid_o                        (valid_o_2_19),
    .ready_i                        (ready_i_2_19)
);


always@(*) begin
    data_i_2_19[3] = data_o_2_18[4];
    valid_i_2_19[3] = valid_o_2_18[4];
    ready_i_2_19[3] = ready_o_2_18[4];
    data_i_2_19[4] = data_o_2_20[3];
    valid_i_2_19[4] = valid_o_2_20[3];
    ready_i_2_19[4] = ready_o_2_20[3];
    data_i_2_19[1] = data_o_1_19[2];
    valid_i_2_19[1] = valid_o_1_19[2];
    ready_i_2_19[1] = ready_o_1_19[2];
    data_i_2_19[2] = data_o_3_19[1];
    valid_i_2_19[2] = valid_o_3_19[1];
    ready_i_2_19[2] = ready_o_3_19[1];
    data_i_2_19[0] = data_i[2][19];
    valid_i_2_19[0] = valid_i[2][19];
    ready_i_2_19[0] = ready_i[2][19];
end


/*Router 2,20*/    
merge_router #(
    .input_mask                     (input_mask_2_20),
    .output_sel                     (output_sel_2_20)
)router202(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_2_20),
    .valid_i                        (valid_i_2_20),
    .ready_o                        (ready_o_2_20),
    .data_o                         (data_o_2_20),
    .valid_o                        (valid_o_2_20),
    .ready_i                        (ready_i_2_20)
);


always@(*) begin
    data_i_2_20[3] = data_o_2_19[4];
    valid_i_2_20[3] = valid_o_2_19[4];
    ready_i_2_20[3] = ready_o_2_19[4];
    data_i_2_20[4] = data_o_2_21[3];
    valid_i_2_20[4] = valid_o_2_21[3];
    ready_i_2_20[4] = ready_o_2_21[3];
    data_i_2_20[1] = data_o_1_20[2];
    valid_i_2_20[1] = valid_o_1_20[2];
    ready_i_2_20[1] = ready_o_1_20[2];
    data_i_2_20[2] = data_o_3_20[1];
    valid_i_2_20[2] = valid_o_3_20[1];
    ready_i_2_20[2] = ready_o_3_20[1];
    data_i_2_20[0] = data_i[2][20];
    valid_i_2_20[0] = valid_i[2][20];
    ready_i_2_20[0] = ready_i[2][20];
end


/*Router 2,21*/    
merge_router #(
    .input_mask                     (input_mask_2_21),
    .output_sel                     (output_sel_2_21)
)router212(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_2_21),
    .valid_i                        (valid_i_2_21),
    .ready_o                        (ready_o_2_21),
    .data_o                         (data_o_2_21),
    .valid_o                        (valid_o_2_21),
    .ready_i                        (ready_i_2_21)
);


always@(*) begin
    data_i_2_21[3] = data_o_2_20[4];
    valid_i_2_21[3] = valid_o_2_20[4];
    ready_i_2_21[3] = ready_o_2_20[4];
    data_i_2_21[4] = data_o_2_22[3];
    valid_i_2_21[4] = valid_o_2_22[3];
    ready_i_2_21[4] = ready_o_2_22[3];
    data_i_2_21[1] = data_o_1_21[2];
    valid_i_2_21[1] = valid_o_1_21[2];
    ready_i_2_21[1] = ready_o_1_21[2];
    data_i_2_21[2] = data_o_3_21[1];
    valid_i_2_21[2] = valid_o_3_21[1];
    ready_i_2_21[2] = ready_o_3_21[1];
    data_i_2_21[0] = data_i[2][21];
    valid_i_2_21[0] = valid_i[2][21];
    ready_i_2_21[0] = ready_i[2][21];
end


/*Router 2,22*/    
merge_router #(
    .input_mask                     (input_mask_2_22),
    .output_sel                     (output_sel_2_22)
)router222(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_2_22),
    .valid_i                        (valid_i_2_22),
    .ready_o                        (ready_o_2_22),
    .data_o                         (data_o_2_22),
    .valid_o                        (valid_o_2_22),
    .ready_i                        (ready_i_2_22)
);


always@(*) begin
    data_i_2_22[3] = data_o_2_21[4];
    valid_i_2_22[3] = valid_o_2_21[4];
    ready_i_2_22[3] = ready_o_2_21[4];
    data_i_2_22[4] = data_o_2_23[3];
    valid_i_2_22[4] = valid_o_2_23[3];
    ready_i_2_22[4] = ready_o_2_23[3];
    data_i_2_22[1] = data_o_1_22[2];
    valid_i_2_22[1] = valid_o_1_22[2];
    ready_i_2_22[1] = ready_o_1_22[2];
    data_i_2_22[2] = data_o_3_22[1];
    valid_i_2_22[2] = valid_o_3_22[1];
    ready_i_2_22[2] = ready_o_3_22[1];
    data_i_2_22[0] = data_i[2][22];
    valid_i_2_22[0] = valid_i[2][22];
    ready_i_2_22[0] = ready_i[2][22];
end


/*Router 2,23*/    
merge_router #(
    .input_mask                     (input_mask_2_23),
    .output_sel                     (output_sel_2_23)
)router232(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_2_23),
    .valid_i                        (valid_i_2_23),
    .ready_o                        (ready_o_2_23),
    .data_o                         (data_o_2_23),
    .valid_o                        (valid_o_2_23),
    .ready_i                        (ready_i_2_23)
);


always@(*) begin
    data_i_2_23[3] = data_o_2_22[4];
    valid_i_2_23[3] = valid_o_2_22[4];
    ready_i_2_23[3] = ready_o_2_22[4];
    data_i_2_23[4] = data_o_2_24[3];
    valid_i_2_23[4] = valid_o_2_24[3];
    ready_i_2_23[4] = ready_o_2_24[3];
    data_i_2_23[1] = data_o_1_23[2];
    valid_i_2_23[1] = valid_o_1_23[2];
    ready_i_2_23[1] = ready_o_1_23[2];
    data_i_2_23[2] = data_o_3_23[1];
    valid_i_2_23[2] = valid_o_3_23[1];
    ready_i_2_23[2] = ready_o_3_23[1];
    data_i_2_23[0] = data_i[2][23];
    valid_i_2_23[0] = valid_i[2][23];
    ready_i_2_23[0] = ready_i[2][23];
end


/*Router 2,24*/    
merge_router #(
    .input_mask                     (input_mask_2_24),
    .output_sel                     (output_sel_2_24)
)router242(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_2_24),
    .valid_i                        (valid_i_2_24),
    .ready_o                        (ready_o_2_24),
    .data_o                         (data_o_2_24),
    .valid_o                        (valid_o_2_24),
    .ready_i                        (ready_i_2_24)
);


always@(*) begin
    data_i_2_24[3] = data_o_2_23[4];
    valid_i_2_24[3] = valid_o_2_23[4];
    ready_i_2_24[3] = ready_o_2_23[4];
    data_i_2_24[1] = data_o_1_24[2];
    valid_i_2_24[1] = valid_o_1_24[2];
    ready_i_2_24[1] = ready_o_1_24[2];
    data_i_2_24[2] = data_o_3_24[1];
    valid_i_2_24[2] = valid_o_3_24[1];
    ready_i_2_24[2] = ready_o_3_24[1];
    data_i_2_24[0] = data_i[2][24];
    valid_i_2_24[0] = valid_i[2][24];
    ready_i_2_24[0] = ready_i[2][24];
end


/*Router 3,0*/    
merge_router #(
    .input_mask                     (input_mask_3_0),
    .output_sel                     (output_sel_3_0)
)router3(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_3_0),
    .valid_i                        (valid_i_3_0),
    .ready_o                        (ready_o_3_0),
    .data_o                         (data_o_3_0),
    .valid_o                        (valid_o_3_0),
    .ready_i                        (ready_i_3_0)
);


always@(*) begin
    data_i_3_0[4] = data_o_3_1[3];
    valid_i_3_0[4] = valid_o_3_1[3];
    ready_i_3_0[4] = ready_o_3_1[3];
    data_i_3_0[1] = data_o_2_0[2];
    valid_i_3_0[1] = valid_o_2_0[2];
    ready_i_3_0[1] = ready_o_2_0[2];
    data_i_3_0[2] = data_o_4_0[1];
    valid_i_3_0[2] = valid_o_4_0[1];
    ready_i_3_0[2] = ready_o_4_0[1];
    data_i_3_0[0] = data_i[3][0];
    valid_i_3_0[0] = valid_i[3][0];
    ready_i_3_0[0] = ready_i[3][0];
end


/*Router 3,1*/    
merge_router #(
    .input_mask                     (input_mask_3_1),
    .output_sel                     (output_sel_3_1)
)router13(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_3_1),
    .valid_i                        (valid_i_3_1),
    .ready_o                        (ready_o_3_1),
    .data_o                         (data_o_3_1),
    .valid_o                        (valid_o_3_1),
    .ready_i                        (ready_i_3_1)
);


always@(*) begin
    data_i_3_1[3] = data_o_3_0[4];
    valid_i_3_1[3] = valid_o_3_0[4];
    ready_i_3_1[3] = ready_o_3_0[4];
    data_i_3_1[4] = data_o_3_2[3];
    valid_i_3_1[4] = valid_o_3_2[3];
    ready_i_3_1[4] = ready_o_3_2[3];
    data_i_3_1[1] = data_o_2_1[2];
    valid_i_3_1[1] = valid_o_2_1[2];
    ready_i_3_1[1] = ready_o_2_1[2];
    data_i_3_1[2] = data_o_4_1[1];
    valid_i_3_1[2] = valid_o_4_1[1];
    ready_i_3_1[2] = ready_o_4_1[1];
    data_i_3_1[0] = data_i[3][1];
    valid_i_3_1[0] = valid_i[3][1];
    ready_i_3_1[0] = ready_i[3][1];
end


/*Router 3,2*/    
merge_router #(
    .input_mask                     (input_mask_3_2),
    .output_sel                     (output_sel_3_2)
)router23(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_3_2),
    .valid_i                        (valid_i_3_2),
    .ready_o                        (ready_o_3_2),
    .data_o                         (data_o_3_2),
    .valid_o                        (valid_o_3_2),
    .ready_i                        (ready_i_3_2)
);


always@(*) begin
    data_i_3_2[3] = data_o_3_1[4];
    valid_i_3_2[3] = valid_o_3_1[4];
    ready_i_3_2[3] = ready_o_3_1[4];
    data_i_3_2[4] = data_o_3_3[3];
    valid_i_3_2[4] = valid_o_3_3[3];
    ready_i_3_2[4] = ready_o_3_3[3];
    data_i_3_2[1] = data_o_2_2[2];
    valid_i_3_2[1] = valid_o_2_2[2];
    ready_i_3_2[1] = ready_o_2_2[2];
    data_i_3_2[2] = data_o_4_2[1];
    valid_i_3_2[2] = valid_o_4_2[1];
    ready_i_3_2[2] = ready_o_4_2[1];
    data_i_3_2[0] = data_i[3][2];
    valid_i_3_2[0] = valid_i[3][2];
    ready_i_3_2[0] = ready_i[3][2];
end


/*Router 3,3*/    
merge_router #(
    .input_mask                     (input_mask_3_3),
    .output_sel                     (output_sel_3_3)
)router33(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_3_3),
    .valid_i                        (valid_i_3_3),
    .ready_o                        (ready_o_3_3),
    .data_o                         (data_o_3_3),
    .valid_o                        (valid_o_3_3),
    .ready_i                        (ready_i_3_3)
);


always@(*) begin
    data_i_3_3[3] = data_o_3_2[4];
    valid_i_3_3[3] = valid_o_3_2[4];
    ready_i_3_3[3] = ready_o_3_2[4];
    data_i_3_3[4] = data_o_3_4[3];
    valid_i_3_3[4] = valid_o_3_4[3];
    ready_i_3_3[4] = ready_o_3_4[3];
    data_i_3_3[1] = data_o_2_3[2];
    valid_i_3_3[1] = valid_o_2_3[2];
    ready_i_3_3[1] = ready_o_2_3[2];
    data_i_3_3[2] = data_o_4_3[1];
    valid_i_3_3[2] = valid_o_4_3[1];
    ready_i_3_3[2] = ready_o_4_3[1];
    data_i_3_3[0] = data_i[3][3];
    valid_i_3_3[0] = valid_i[3][3];
    ready_i_3_3[0] = ready_i[3][3];
end


/*Router 3,4*/    
merge_router #(
    .input_mask                     (input_mask_3_4),
    .output_sel                     (output_sel_3_4)
)router43(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_3_4),
    .valid_i                        (valid_i_3_4),
    .ready_o                        (ready_o_3_4),
    .data_o                         (data_o_3_4),
    .valid_o                        (valid_o_3_4),
    .ready_i                        (ready_i_3_4)
);


always@(*) begin
    data_i_3_4[3] = data_o_3_3[4];
    valid_i_3_4[3] = valid_o_3_3[4];
    ready_i_3_4[3] = ready_o_3_3[4];
    data_i_3_4[4] = data_o_3_5[3];
    valid_i_3_4[4] = valid_o_3_5[3];
    ready_i_3_4[4] = ready_o_3_5[3];
    data_i_3_4[1] = data_o_2_4[2];
    valid_i_3_4[1] = valid_o_2_4[2];
    ready_i_3_4[1] = ready_o_2_4[2];
    data_i_3_4[2] = data_o_4_4[1];
    valid_i_3_4[2] = valid_o_4_4[1];
    ready_i_3_4[2] = ready_o_4_4[1];
    data_i_3_4[0] = data_i[3][4];
    valid_i_3_4[0] = valid_i[3][4];
    ready_i_3_4[0] = ready_i[3][4];
end


/*Router 3,5*/    
merge_router #(
    .input_mask                     (input_mask_3_5),
    .output_sel                     (output_sel_3_5)
)router53(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_3_5),
    .valid_i                        (valid_i_3_5),
    .ready_o                        (ready_o_3_5),
    .data_o                         (data_o_3_5),
    .valid_o                        (valid_o_3_5),
    .ready_i                        (ready_i_3_5)
);


always@(*) begin
    data_i_3_5[3] = data_o_3_4[4];
    valid_i_3_5[3] = valid_o_3_4[4];
    ready_i_3_5[3] = ready_o_3_4[4];
    data_i_3_5[4] = data_o_3_6[3];
    valid_i_3_5[4] = valid_o_3_6[3];
    ready_i_3_5[4] = ready_o_3_6[3];
    data_i_3_5[1] = data_o_2_5[2];
    valid_i_3_5[1] = valid_o_2_5[2];
    ready_i_3_5[1] = ready_o_2_5[2];
    data_i_3_5[2] = data_o_4_5[1];
    valid_i_3_5[2] = valid_o_4_5[1];
    ready_i_3_5[2] = ready_o_4_5[1];
    data_i_3_5[0] = data_i[3][5];
    valid_i_3_5[0] = valid_i[3][5];
    ready_i_3_5[0] = ready_i[3][5];
end


/*Router 3,6*/    
merge_router #(
    .input_mask                     (input_mask_3_6),
    .output_sel                     (output_sel_3_6)
)router63(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_3_6),
    .valid_i                        (valid_i_3_6),
    .ready_o                        (ready_o_3_6),
    .data_o                         (data_o_3_6),
    .valid_o                        (valid_o_3_6),
    .ready_i                        (ready_i_3_6)
);


always@(*) begin
    data_i_3_6[3] = data_o_3_5[4];
    valid_i_3_6[3] = valid_o_3_5[4];
    ready_i_3_6[3] = ready_o_3_5[4];
    data_i_3_6[4] = data_o_3_7[3];
    valid_i_3_6[4] = valid_o_3_7[3];
    ready_i_3_6[4] = ready_o_3_7[3];
    data_i_3_6[1] = data_o_2_6[2];
    valid_i_3_6[1] = valid_o_2_6[2];
    ready_i_3_6[1] = ready_o_2_6[2];
    data_i_3_6[2] = data_o_4_6[1];
    valid_i_3_6[2] = valid_o_4_6[1];
    ready_i_3_6[2] = ready_o_4_6[1];
    data_i_3_6[0] = data_i[3][6];
    valid_i_3_6[0] = valid_i[3][6];
    ready_i_3_6[0] = ready_i[3][6];
end


/*Router 3,7*/    
merge_router #(
    .input_mask                     (input_mask_3_7),
    .output_sel                     (output_sel_3_7)
)router73(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_3_7),
    .valid_i                        (valid_i_3_7),
    .ready_o                        (ready_o_3_7),
    .data_o                         (data_o_3_7),
    .valid_o                        (valid_o_3_7),
    .ready_i                        (ready_i_3_7)
);


always@(*) begin
    data_i_3_7[3] = data_o_3_6[4];
    valid_i_3_7[3] = valid_o_3_6[4];
    ready_i_3_7[3] = ready_o_3_6[4];
    data_i_3_7[4] = data_o_3_8[3];
    valid_i_3_7[4] = valid_o_3_8[3];
    ready_i_3_7[4] = ready_o_3_8[3];
    data_i_3_7[1] = data_o_2_7[2];
    valid_i_3_7[1] = valid_o_2_7[2];
    ready_i_3_7[1] = ready_o_2_7[2];
    data_i_3_7[2] = data_o_4_7[1];
    valid_i_3_7[2] = valid_o_4_7[1];
    ready_i_3_7[2] = ready_o_4_7[1];
    data_i_3_7[0] = data_i[3][7];
    valid_i_3_7[0] = valid_i[3][7];
    ready_i_3_7[0] = ready_i[3][7];
end


/*Router 3,8*/    
merge_router #(
    .input_mask                     (input_mask_3_8),
    .output_sel                     (output_sel_3_8)
)router83(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_3_8),
    .valid_i                        (valid_i_3_8),
    .ready_o                        (ready_o_3_8),
    .data_o                         (data_o_3_8),
    .valid_o                        (valid_o_3_8),
    .ready_i                        (ready_i_3_8)
);


always@(*) begin
    data_i_3_8[3] = data_o_3_7[4];
    valid_i_3_8[3] = valid_o_3_7[4];
    ready_i_3_8[3] = ready_o_3_7[4];
    data_i_3_8[4] = data_o_3_9[3];
    valid_i_3_8[4] = valid_o_3_9[3];
    ready_i_3_8[4] = ready_o_3_9[3];
    data_i_3_8[1] = data_o_2_8[2];
    valid_i_3_8[1] = valid_o_2_8[2];
    ready_i_3_8[1] = ready_o_2_8[2];
    data_i_3_8[2] = data_o_4_8[1];
    valid_i_3_8[2] = valid_o_4_8[1];
    ready_i_3_8[2] = ready_o_4_8[1];
    data_i_3_8[0] = data_i[3][8];
    valid_i_3_8[0] = valid_i[3][8];
    ready_i_3_8[0] = ready_i[3][8];
end


/*Router 3,9*/    
merge_router #(
    .input_mask                     (input_mask_3_9),
    .output_sel                     (output_sel_3_9)
)router93(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_3_9),
    .valid_i                        (valid_i_3_9),
    .ready_o                        (ready_o_3_9),
    .data_o                         (data_o_3_9),
    .valid_o                        (valid_o_3_9),
    .ready_i                        (ready_i_3_9)
);


always@(*) begin
    data_i_3_9[3] = data_o_3_8[4];
    valid_i_3_9[3] = valid_o_3_8[4];
    ready_i_3_9[3] = ready_o_3_8[4];
    data_i_3_9[4] = data_o_3_10[3];
    valid_i_3_9[4] = valid_o_3_10[3];
    ready_i_3_9[4] = ready_o_3_10[3];
    data_i_3_9[1] = data_o_2_9[2];
    valid_i_3_9[1] = valid_o_2_9[2];
    ready_i_3_9[1] = ready_o_2_9[2];
    data_i_3_9[2] = data_o_4_9[1];
    valid_i_3_9[2] = valid_o_4_9[1];
    ready_i_3_9[2] = ready_o_4_9[1];
    data_i_3_9[0] = data_i[3][9];
    valid_i_3_9[0] = valid_i[3][9];
    ready_i_3_9[0] = ready_i[3][9];
end


/*Router 3,10*/    
merge_router #(
    .input_mask                     (input_mask_3_10),
    .output_sel                     (output_sel_3_10)
)router103(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_3_10),
    .valid_i                        (valid_i_3_10),
    .ready_o                        (ready_o_3_10),
    .data_o                         (data_o_3_10),
    .valid_o                        (valid_o_3_10),
    .ready_i                        (ready_i_3_10)
);


always@(*) begin
    data_i_3_10[3] = data_o_3_9[4];
    valid_i_3_10[3] = valid_o_3_9[4];
    ready_i_3_10[3] = ready_o_3_9[4];
    data_i_3_10[4] = data_o_3_11[3];
    valid_i_3_10[4] = valid_o_3_11[3];
    ready_i_3_10[4] = ready_o_3_11[3];
    data_i_3_10[1] = data_o_2_10[2];
    valid_i_3_10[1] = valid_o_2_10[2];
    ready_i_3_10[1] = ready_o_2_10[2];
    data_i_3_10[2] = data_o_4_10[1];
    valid_i_3_10[2] = valid_o_4_10[1];
    ready_i_3_10[2] = ready_o_4_10[1];
    data_i_3_10[0] = data_i[3][10];
    valid_i_3_10[0] = valid_i[3][10];
    ready_i_3_10[0] = ready_i[3][10];
end


/*Router 3,11*/    
merge_router #(
    .input_mask                     (input_mask_3_11),
    .output_sel                     (output_sel_3_11)
)router113(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_3_11),
    .valid_i                        (valid_i_3_11),
    .ready_o                        (ready_o_3_11),
    .data_o                         (data_o_3_11),
    .valid_o                        (valid_o_3_11),
    .ready_i                        (ready_i_3_11)
);


always@(*) begin
    data_i_3_11[3] = data_o_3_10[4];
    valid_i_3_11[3] = valid_o_3_10[4];
    ready_i_3_11[3] = ready_o_3_10[4];
    data_i_3_11[4] = data_o_3_12[3];
    valid_i_3_11[4] = valid_o_3_12[3];
    ready_i_3_11[4] = ready_o_3_12[3];
    data_i_3_11[1] = data_o_2_11[2];
    valid_i_3_11[1] = valid_o_2_11[2];
    ready_i_3_11[1] = ready_o_2_11[2];
    data_i_3_11[2] = data_o_4_11[1];
    valid_i_3_11[2] = valid_o_4_11[1];
    ready_i_3_11[2] = ready_o_4_11[1];
    data_i_3_11[0] = data_i[3][11];
    valid_i_3_11[0] = valid_i[3][11];
    ready_i_3_11[0] = ready_i[3][11];
end


/*Router 3,12*/    
merge_router #(
    .input_mask                     (input_mask_3_12),
    .output_sel                     (output_sel_3_12)
)router123(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_3_12),
    .valid_i                        (valid_i_3_12),
    .ready_o                        (ready_o_3_12),
    .data_o                         (data_o_3_12),
    .valid_o                        (valid_o_3_12),
    .ready_i                        (ready_i_3_12)
);


always@(*) begin
    data_i_3_12[3] = data_o_3_11[4];
    valid_i_3_12[3] = valid_o_3_11[4];
    ready_i_3_12[3] = ready_o_3_11[4];
    data_i_3_12[4] = data_o_3_13[3];
    valid_i_3_12[4] = valid_o_3_13[3];
    ready_i_3_12[4] = ready_o_3_13[3];
    data_i_3_12[1] = data_o_2_12[2];
    valid_i_3_12[1] = valid_o_2_12[2];
    ready_i_3_12[1] = ready_o_2_12[2];
    data_i_3_12[2] = data_o_4_12[1];
    valid_i_3_12[2] = valid_o_4_12[1];
    ready_i_3_12[2] = ready_o_4_12[1];
    data_i_3_12[0] = data_i[3][12];
    valid_i_3_12[0] = valid_i[3][12];
    ready_i_3_12[0] = ready_i[3][12];
end


/*Router 3,13*/    
merge_router #(
    .input_mask                     (input_mask_3_13),
    .output_sel                     (output_sel_3_13)
)router133(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_3_13),
    .valid_i                        (valid_i_3_13),
    .ready_o                        (ready_o_3_13),
    .data_o                         (data_o_3_13),
    .valid_o                        (valid_o_3_13),
    .ready_i                        (ready_i_3_13)
);


always@(*) begin
    data_i_3_13[3] = data_o_3_12[4];
    valid_i_3_13[3] = valid_o_3_12[4];
    ready_i_3_13[3] = ready_o_3_12[4];
    data_i_3_13[4] = data_o_3_14[3];
    valid_i_3_13[4] = valid_o_3_14[3];
    ready_i_3_13[4] = ready_o_3_14[3];
    data_i_3_13[1] = data_o_2_13[2];
    valid_i_3_13[1] = valid_o_2_13[2];
    ready_i_3_13[1] = ready_o_2_13[2];
    data_i_3_13[2] = data_o_4_13[1];
    valid_i_3_13[2] = valid_o_4_13[1];
    ready_i_3_13[2] = ready_o_4_13[1];
    data_i_3_13[0] = data_i[3][13];
    valid_i_3_13[0] = valid_i[3][13];
    ready_i_3_13[0] = ready_i[3][13];
end


/*Router 3,14*/    
merge_router #(
    .input_mask                     (input_mask_3_14),
    .output_sel                     (output_sel_3_14)
)router143(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_3_14),
    .valid_i                        (valid_i_3_14),
    .ready_o                        (ready_o_3_14),
    .data_o                         (data_o_3_14),
    .valid_o                        (valid_o_3_14),
    .ready_i                        (ready_i_3_14)
);


always@(*) begin
    data_i_3_14[3] = data_o_3_13[4];
    valid_i_3_14[3] = valid_o_3_13[4];
    ready_i_3_14[3] = ready_o_3_13[4];
    data_i_3_14[4] = data_o_3_15[3];
    valid_i_3_14[4] = valid_o_3_15[3];
    ready_i_3_14[4] = ready_o_3_15[3];
    data_i_3_14[1] = data_o_2_14[2];
    valid_i_3_14[1] = valid_o_2_14[2];
    ready_i_3_14[1] = ready_o_2_14[2];
    data_i_3_14[2] = data_o_4_14[1];
    valid_i_3_14[2] = valid_o_4_14[1];
    ready_i_3_14[2] = ready_o_4_14[1];
    data_i_3_14[0] = data_i[3][14];
    valid_i_3_14[0] = valid_i[3][14];
    ready_i_3_14[0] = ready_i[3][14];
end


/*Router 3,15*/    
merge_router #(
    .input_mask                     (input_mask_3_15),
    .output_sel                     (output_sel_3_15)
)router153(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_3_15),
    .valid_i                        (valid_i_3_15),
    .ready_o                        (ready_o_3_15),
    .data_o                         (data_o_3_15),
    .valid_o                        (valid_o_3_15),
    .ready_i                        (ready_i_3_15)
);


always@(*) begin
    data_i_3_15[3] = data_o_3_14[4];
    valid_i_3_15[3] = valid_o_3_14[4];
    ready_i_3_15[3] = ready_o_3_14[4];
    data_i_3_15[4] = data_o_3_16[3];
    valid_i_3_15[4] = valid_o_3_16[3];
    ready_i_3_15[4] = ready_o_3_16[3];
    data_i_3_15[1] = data_o_2_15[2];
    valid_i_3_15[1] = valid_o_2_15[2];
    ready_i_3_15[1] = ready_o_2_15[2];
    data_i_3_15[2] = data_o_4_15[1];
    valid_i_3_15[2] = valid_o_4_15[1];
    ready_i_3_15[2] = ready_o_4_15[1];
    data_i_3_15[0] = data_i[3][15];
    valid_i_3_15[0] = valid_i[3][15];
    ready_i_3_15[0] = ready_i[3][15];
end


/*Router 3,16*/    
merge_router #(
    .input_mask                     (input_mask_3_16),
    .output_sel                     (output_sel_3_16)
)router163(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_3_16),
    .valid_i                        (valid_i_3_16),
    .ready_o                        (ready_o_3_16),
    .data_o                         (data_o_3_16),
    .valid_o                        (valid_o_3_16),
    .ready_i                        (ready_i_3_16)
);


always@(*) begin
    data_i_3_16[3] = data_o_3_15[4];
    valid_i_3_16[3] = valid_o_3_15[4];
    ready_i_3_16[3] = ready_o_3_15[4];
    data_i_3_16[4] = data_o_3_17[3];
    valid_i_3_16[4] = valid_o_3_17[3];
    ready_i_3_16[4] = ready_o_3_17[3];
    data_i_3_16[1] = data_o_2_16[2];
    valid_i_3_16[1] = valid_o_2_16[2];
    ready_i_3_16[1] = ready_o_2_16[2];
    data_i_3_16[2] = data_o_4_16[1];
    valid_i_3_16[2] = valid_o_4_16[1];
    ready_i_3_16[2] = ready_o_4_16[1];
    data_i_3_16[0] = data_i[3][16];
    valid_i_3_16[0] = valid_i[3][16];
    ready_i_3_16[0] = ready_i[3][16];
end


/*Router 3,17*/    
merge_router #(
    .input_mask                     (input_mask_3_17),
    .output_sel                     (output_sel_3_17)
)router173(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_3_17),
    .valid_i                        (valid_i_3_17),
    .ready_o                        (ready_o_3_17),
    .data_o                         (data_o_3_17),
    .valid_o                        (valid_o_3_17),
    .ready_i                        (ready_i_3_17)
);


always@(*) begin
    data_i_3_17[3] = data_o_3_16[4];
    valid_i_3_17[3] = valid_o_3_16[4];
    ready_i_3_17[3] = ready_o_3_16[4];
    data_i_3_17[4] = data_o_3_18[3];
    valid_i_3_17[4] = valid_o_3_18[3];
    ready_i_3_17[4] = ready_o_3_18[3];
    data_i_3_17[1] = data_o_2_17[2];
    valid_i_3_17[1] = valid_o_2_17[2];
    ready_i_3_17[1] = ready_o_2_17[2];
    data_i_3_17[2] = data_o_4_17[1];
    valid_i_3_17[2] = valid_o_4_17[1];
    ready_i_3_17[2] = ready_o_4_17[1];
    data_i_3_17[0] = data_i[3][17];
    valid_i_3_17[0] = valid_i[3][17];
    ready_i_3_17[0] = ready_i[3][17];
end


/*Router 3,18*/    
merge_router #(
    .input_mask                     (input_mask_3_18),
    .output_sel                     (output_sel_3_18)
)router183(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_3_18),
    .valid_i                        (valid_i_3_18),
    .ready_o                        (ready_o_3_18),
    .data_o                         (data_o_3_18),
    .valid_o                        (valid_o_3_18),
    .ready_i                        (ready_i_3_18)
);


always@(*) begin
    data_i_3_18[3] = data_o_3_17[4];
    valid_i_3_18[3] = valid_o_3_17[4];
    ready_i_3_18[3] = ready_o_3_17[4];
    data_i_3_18[4] = data_o_3_19[3];
    valid_i_3_18[4] = valid_o_3_19[3];
    ready_i_3_18[4] = ready_o_3_19[3];
    data_i_3_18[1] = data_o_2_18[2];
    valid_i_3_18[1] = valid_o_2_18[2];
    ready_i_3_18[1] = ready_o_2_18[2];
    data_i_3_18[2] = data_o_4_18[1];
    valid_i_3_18[2] = valid_o_4_18[1];
    ready_i_3_18[2] = ready_o_4_18[1];
    data_i_3_18[0] = data_i[3][18];
    valid_i_3_18[0] = valid_i[3][18];
    ready_i_3_18[0] = ready_i[3][18];
end


/*Router 3,19*/    
merge_router #(
    .input_mask                     (input_mask_3_19),
    .output_sel                     (output_sel_3_19)
)router193(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_3_19),
    .valid_i                        (valid_i_3_19),
    .ready_o                        (ready_o_3_19),
    .data_o                         (data_o_3_19),
    .valid_o                        (valid_o_3_19),
    .ready_i                        (ready_i_3_19)
);


always@(*) begin
    data_i_3_19[3] = data_o_3_18[4];
    valid_i_3_19[3] = valid_o_3_18[4];
    ready_i_3_19[3] = ready_o_3_18[4];
    data_i_3_19[4] = data_o_3_20[3];
    valid_i_3_19[4] = valid_o_3_20[3];
    ready_i_3_19[4] = ready_o_3_20[3];
    data_i_3_19[1] = data_o_2_19[2];
    valid_i_3_19[1] = valid_o_2_19[2];
    ready_i_3_19[1] = ready_o_2_19[2];
    data_i_3_19[2] = data_o_4_19[1];
    valid_i_3_19[2] = valid_o_4_19[1];
    ready_i_3_19[2] = ready_o_4_19[1];
    data_i_3_19[0] = data_i[3][19];
    valid_i_3_19[0] = valid_i[3][19];
    ready_i_3_19[0] = ready_i[3][19];
end


/*Router 3,20*/    
merge_router #(
    .input_mask                     (input_mask_3_20),
    .output_sel                     (output_sel_3_20)
)router203(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_3_20),
    .valid_i                        (valid_i_3_20),
    .ready_o                        (ready_o_3_20),
    .data_o                         (data_o_3_20),
    .valid_o                        (valid_o_3_20),
    .ready_i                        (ready_i_3_20)
);


always@(*) begin
    data_i_3_20[3] = data_o_3_19[4];
    valid_i_3_20[3] = valid_o_3_19[4];
    ready_i_3_20[3] = ready_o_3_19[4];
    data_i_3_20[4] = data_o_3_21[3];
    valid_i_3_20[4] = valid_o_3_21[3];
    ready_i_3_20[4] = ready_o_3_21[3];
    data_i_3_20[1] = data_o_2_20[2];
    valid_i_3_20[1] = valid_o_2_20[2];
    ready_i_3_20[1] = ready_o_2_20[2];
    data_i_3_20[2] = data_o_4_20[1];
    valid_i_3_20[2] = valid_o_4_20[1];
    ready_i_3_20[2] = ready_o_4_20[1];
    data_i_3_20[0] = data_i[3][20];
    valid_i_3_20[0] = valid_i[3][20];
    ready_i_3_20[0] = ready_i[3][20];
end


/*Router 3,21*/    
merge_router #(
    .input_mask                     (input_mask_3_21),
    .output_sel                     (output_sel_3_21)
)router213(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_3_21),
    .valid_i                        (valid_i_3_21),
    .ready_o                        (ready_o_3_21),
    .data_o                         (data_o_3_21),
    .valid_o                        (valid_o_3_21),
    .ready_i                        (ready_i_3_21)
);


always@(*) begin
    data_i_3_21[3] = data_o_3_20[4];
    valid_i_3_21[3] = valid_o_3_20[4];
    ready_i_3_21[3] = ready_o_3_20[4];
    data_i_3_21[4] = data_o_3_22[3];
    valid_i_3_21[4] = valid_o_3_22[3];
    ready_i_3_21[4] = ready_o_3_22[3];
    data_i_3_21[1] = data_o_2_21[2];
    valid_i_3_21[1] = valid_o_2_21[2];
    ready_i_3_21[1] = ready_o_2_21[2];
    data_i_3_21[2] = data_o_4_21[1];
    valid_i_3_21[2] = valid_o_4_21[1];
    ready_i_3_21[2] = ready_o_4_21[1];
    data_i_3_21[0] = data_i[3][21];
    valid_i_3_21[0] = valid_i[3][21];
    ready_i_3_21[0] = ready_i[3][21];
end


/*Router 3,22*/    
merge_router #(
    .input_mask                     (input_mask_3_22),
    .output_sel                     (output_sel_3_22)
)router223(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_3_22),
    .valid_i                        (valid_i_3_22),
    .ready_o                        (ready_o_3_22),
    .data_o                         (data_o_3_22),
    .valid_o                        (valid_o_3_22),
    .ready_i                        (ready_i_3_22)
);


always@(*) begin
    data_i_3_22[3] = data_o_3_21[4];
    valid_i_3_22[3] = valid_o_3_21[4];
    ready_i_3_22[3] = ready_o_3_21[4];
    data_i_3_22[4] = data_o_3_23[3];
    valid_i_3_22[4] = valid_o_3_23[3];
    ready_i_3_22[4] = ready_o_3_23[3];
    data_i_3_22[1] = data_o_2_22[2];
    valid_i_3_22[1] = valid_o_2_22[2];
    ready_i_3_22[1] = ready_o_2_22[2];
    data_i_3_22[2] = data_o_4_22[1];
    valid_i_3_22[2] = valid_o_4_22[1];
    ready_i_3_22[2] = ready_o_4_22[1];
    data_i_3_22[0] = data_i[3][22];
    valid_i_3_22[0] = valid_i[3][22];
    ready_i_3_22[0] = ready_i[3][22];
end


/*Router 3,23*/    
merge_router #(
    .input_mask                     (input_mask_3_23),
    .output_sel                     (output_sel_3_23)
)router233(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_3_23),
    .valid_i                        (valid_i_3_23),
    .ready_o                        (ready_o_3_23),
    .data_o                         (data_o_3_23),
    .valid_o                        (valid_o_3_23),
    .ready_i                        (ready_i_3_23)
);


always@(*) begin
    data_i_3_23[3] = data_o_3_22[4];
    valid_i_3_23[3] = valid_o_3_22[4];
    ready_i_3_23[3] = ready_o_3_22[4];
    data_i_3_23[4] = data_o_3_24[3];
    valid_i_3_23[4] = valid_o_3_24[3];
    ready_i_3_23[4] = ready_o_3_24[3];
    data_i_3_23[1] = data_o_2_23[2];
    valid_i_3_23[1] = valid_o_2_23[2];
    ready_i_3_23[1] = ready_o_2_23[2];
    data_i_3_23[2] = data_o_4_23[1];
    valid_i_3_23[2] = valid_o_4_23[1];
    ready_i_3_23[2] = ready_o_4_23[1];
    data_i_3_23[0] = data_i[3][23];
    valid_i_3_23[0] = valid_i[3][23];
    ready_i_3_23[0] = ready_i[3][23];
end


/*Router 3,24*/    
merge_router #(
    .input_mask                     (input_mask_3_24),
    .output_sel                     (output_sel_3_24)
)router243(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_3_24),
    .valid_i                        (valid_i_3_24),
    .ready_o                        (ready_o_3_24),
    .data_o                         (data_o_3_24),
    .valid_o                        (valid_o_3_24),
    .ready_i                        (ready_i_3_24)
);


always@(*) begin
    data_i_3_24[3] = data_o_3_23[4];
    valid_i_3_24[3] = valid_o_3_23[4];
    ready_i_3_24[3] = ready_o_3_23[4];
    data_i_3_24[1] = data_o_2_24[2];
    valid_i_3_24[1] = valid_o_2_24[2];
    ready_i_3_24[1] = ready_o_2_24[2];
    data_i_3_24[2] = data_o_4_24[1];
    valid_i_3_24[2] = valid_o_4_24[1];
    ready_i_3_24[2] = ready_o_4_24[1];
    data_i_3_24[0] = data_i[3][24];
    valid_i_3_24[0] = valid_i[3][24];
    ready_i_3_24[0] = ready_i[3][24];
end


/*Router 4,0*/    
merge_router #(
    .input_mask                     (input_mask_4_0),
    .output_sel                     (output_sel_4_0)
)router4(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_4_0),
    .valid_i                        (valid_i_4_0),
    .ready_o                        (ready_o_4_0),
    .data_o                         (data_o_4_0),
    .valid_o                        (valid_o_4_0),
    .ready_i                        (ready_i_4_0)
);


always@(*) begin
    data_i_4_0[4] = data_o_4_1[3];
    valid_i_4_0[4] = valid_o_4_1[3];
    ready_i_4_0[4] = ready_o_4_1[3];
    data_i_4_0[1] = data_o_3_0[2];
    valid_i_4_0[1] = valid_o_3_0[2];
    ready_i_4_0[1] = ready_o_3_0[2];
    data_i_4_0[2] = data_o_5_0[1];
    valid_i_4_0[2] = valid_o_5_0[1];
    ready_i_4_0[2] = ready_o_5_0[1];
    data_i_4_0[0] = data_i[4][0];
    valid_i_4_0[0] = valid_i[4][0];
    ready_i_4_0[0] = ready_i[4][0];
end


/*Router 4,1*/    
merge_router #(
    .input_mask                     (input_mask_4_1),
    .output_sel                     (output_sel_4_1)
)router14(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_4_1),
    .valid_i                        (valid_i_4_1),
    .ready_o                        (ready_o_4_1),
    .data_o                         (data_o_4_1),
    .valid_o                        (valid_o_4_1),
    .ready_i                        (ready_i_4_1)
);


always@(*) begin
    data_i_4_1[3] = data_o_4_0[4];
    valid_i_4_1[3] = valid_o_4_0[4];
    ready_i_4_1[3] = ready_o_4_0[4];
    data_i_4_1[4] = data_o_4_2[3];
    valid_i_4_1[4] = valid_o_4_2[3];
    ready_i_4_1[4] = ready_o_4_2[3];
    data_i_4_1[1] = data_o_3_1[2];
    valid_i_4_1[1] = valid_o_3_1[2];
    ready_i_4_1[1] = ready_o_3_1[2];
    data_i_4_1[2] = data_o_5_1[1];
    valid_i_4_1[2] = valid_o_5_1[1];
    ready_i_4_1[2] = ready_o_5_1[1];
    data_i_4_1[0] = data_i[4][1];
    valid_i_4_1[0] = valid_i[4][1];
    ready_i_4_1[0] = ready_i[4][1];
end


/*Router 4,2*/    
merge_router #(
    .input_mask                     (input_mask_4_2),
    .output_sel                     (output_sel_4_2)
)router24(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_4_2),
    .valid_i                        (valid_i_4_2),
    .ready_o                        (ready_o_4_2),
    .data_o                         (data_o_4_2),
    .valid_o                        (valid_o_4_2),
    .ready_i                        (ready_i_4_2)
);


always@(*) begin
    data_i_4_2[3] = data_o_4_1[4];
    valid_i_4_2[3] = valid_o_4_1[4];
    ready_i_4_2[3] = ready_o_4_1[4];
    data_i_4_2[4] = data_o_4_3[3];
    valid_i_4_2[4] = valid_o_4_3[3];
    ready_i_4_2[4] = ready_o_4_3[3];
    data_i_4_2[1] = data_o_3_2[2];
    valid_i_4_2[1] = valid_o_3_2[2];
    ready_i_4_2[1] = ready_o_3_2[2];
    data_i_4_2[2] = data_o_5_2[1];
    valid_i_4_2[2] = valid_o_5_2[1];
    ready_i_4_2[2] = ready_o_5_2[1];
    data_i_4_2[0] = data_i[4][2];
    valid_i_4_2[0] = valid_i[4][2];
    ready_i_4_2[0] = ready_i[4][2];
end


/*Router 4,3*/    
merge_router #(
    .input_mask                     (input_mask_4_3),
    .output_sel                     (output_sel_4_3)
)router34(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_4_3),
    .valid_i                        (valid_i_4_3),
    .ready_o                        (ready_o_4_3),
    .data_o                         (data_o_4_3),
    .valid_o                        (valid_o_4_3),
    .ready_i                        (ready_i_4_3)
);


always@(*) begin
    data_i_4_3[3] = data_o_4_2[4];
    valid_i_4_3[3] = valid_o_4_2[4];
    ready_i_4_3[3] = ready_o_4_2[4];
    data_i_4_3[4] = data_o_4_4[3];
    valid_i_4_3[4] = valid_o_4_4[3];
    ready_i_4_3[4] = ready_o_4_4[3];
    data_i_4_3[1] = data_o_3_3[2];
    valid_i_4_3[1] = valid_o_3_3[2];
    ready_i_4_3[1] = ready_o_3_3[2];
    data_i_4_3[2] = data_o_5_3[1];
    valid_i_4_3[2] = valid_o_5_3[1];
    ready_i_4_3[2] = ready_o_5_3[1];
    data_i_4_3[0] = data_i[4][3];
    valid_i_4_3[0] = valid_i[4][3];
    ready_i_4_3[0] = ready_i[4][3];
end


/*Router 4,4*/    
merge_router #(
    .input_mask                     (input_mask_4_4),
    .output_sel                     (output_sel_4_4)
)router44(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_4_4),
    .valid_i                        (valid_i_4_4),
    .ready_o                        (ready_o_4_4),
    .data_o                         (data_o_4_4),
    .valid_o                        (valid_o_4_4),
    .ready_i                        (ready_i_4_4)
);


always@(*) begin
    data_i_4_4[3] = data_o_4_3[4];
    valid_i_4_4[3] = valid_o_4_3[4];
    ready_i_4_4[3] = ready_o_4_3[4];
    data_i_4_4[4] = data_o_4_5[3];
    valid_i_4_4[4] = valid_o_4_5[3];
    ready_i_4_4[4] = ready_o_4_5[3];
    data_i_4_4[1] = data_o_3_4[2];
    valid_i_4_4[1] = valid_o_3_4[2];
    ready_i_4_4[1] = ready_o_3_4[2];
    data_i_4_4[2] = data_o_5_4[1];
    valid_i_4_4[2] = valid_o_5_4[1];
    ready_i_4_4[2] = ready_o_5_4[1];
    data_i_4_4[0] = data_i[4][4];
    valid_i_4_4[0] = valid_i[4][4];
    ready_i_4_4[0] = ready_i[4][4];
end


/*Router 4,5*/    
merge_router #(
    .input_mask                     (input_mask_4_5),
    .output_sel                     (output_sel_4_5)
)router54(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_4_5),
    .valid_i                        (valid_i_4_5),
    .ready_o                        (ready_o_4_5),
    .data_o                         (data_o_4_5),
    .valid_o                        (valid_o_4_5),
    .ready_i                        (ready_i_4_5)
);


always@(*) begin
    data_i_4_5[3] = data_o_4_4[4];
    valid_i_4_5[3] = valid_o_4_4[4];
    ready_i_4_5[3] = ready_o_4_4[4];
    data_i_4_5[4] = data_o_4_6[3];
    valid_i_4_5[4] = valid_o_4_6[3];
    ready_i_4_5[4] = ready_o_4_6[3];
    data_i_4_5[1] = data_o_3_5[2];
    valid_i_4_5[1] = valid_o_3_5[2];
    ready_i_4_5[1] = ready_o_3_5[2];
    data_i_4_5[2] = data_o_5_5[1];
    valid_i_4_5[2] = valid_o_5_5[1];
    ready_i_4_5[2] = ready_o_5_5[1];
    data_i_4_5[0] = data_i[4][5];
    valid_i_4_5[0] = valid_i[4][5];
    ready_i_4_5[0] = ready_i[4][5];
end


/*Router 4,6*/    
merge_router #(
    .input_mask                     (input_mask_4_6),
    .output_sel                     (output_sel_4_6)
)router64(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_4_6),
    .valid_i                        (valid_i_4_6),
    .ready_o                        (ready_o_4_6),
    .data_o                         (data_o_4_6),
    .valid_o                        (valid_o_4_6),
    .ready_i                        (ready_i_4_6)
);


always@(*) begin
    data_i_4_6[3] = data_o_4_5[4];
    valid_i_4_6[3] = valid_o_4_5[4];
    ready_i_4_6[3] = ready_o_4_5[4];
    data_i_4_6[4] = data_o_4_7[3];
    valid_i_4_6[4] = valid_o_4_7[3];
    ready_i_4_6[4] = ready_o_4_7[3];
    data_i_4_6[1] = data_o_3_6[2];
    valid_i_4_6[1] = valid_o_3_6[2];
    ready_i_4_6[1] = ready_o_3_6[2];
    data_i_4_6[2] = data_o_5_6[1];
    valid_i_4_6[2] = valid_o_5_6[1];
    ready_i_4_6[2] = ready_o_5_6[1];
    data_i_4_6[0] = data_i[4][6];
    valid_i_4_6[0] = valid_i[4][6];
    ready_i_4_6[0] = ready_i[4][6];
end


/*Router 4,7*/    
merge_router #(
    .input_mask                     (input_mask_4_7),
    .output_sel                     (output_sel_4_7)
)router74(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_4_7),
    .valid_i                        (valid_i_4_7),
    .ready_o                        (ready_o_4_7),
    .data_o                         (data_o_4_7),
    .valid_o                        (valid_o_4_7),
    .ready_i                        (ready_i_4_7)
);


always@(*) begin
    data_i_4_7[3] = data_o_4_6[4];
    valid_i_4_7[3] = valid_o_4_6[4];
    ready_i_4_7[3] = ready_o_4_6[4];
    data_i_4_7[4] = data_o_4_8[3];
    valid_i_4_7[4] = valid_o_4_8[3];
    ready_i_4_7[4] = ready_o_4_8[3];
    data_i_4_7[1] = data_o_3_7[2];
    valid_i_4_7[1] = valid_o_3_7[2];
    ready_i_4_7[1] = ready_o_3_7[2];
    data_i_4_7[2] = data_o_5_7[1];
    valid_i_4_7[2] = valid_o_5_7[1];
    ready_i_4_7[2] = ready_o_5_7[1];
    data_i_4_7[0] = data_i[4][7];
    valid_i_4_7[0] = valid_i[4][7];
    ready_i_4_7[0] = ready_i[4][7];
end


/*Router 4,8*/    
merge_router #(
    .input_mask                     (input_mask_4_8),
    .output_sel                     (output_sel_4_8)
)router84(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_4_8),
    .valid_i                        (valid_i_4_8),
    .ready_o                        (ready_o_4_8),
    .data_o                         (data_o_4_8),
    .valid_o                        (valid_o_4_8),
    .ready_i                        (ready_i_4_8)
);


always@(*) begin
    data_i_4_8[3] = data_o_4_7[4];
    valid_i_4_8[3] = valid_o_4_7[4];
    ready_i_4_8[3] = ready_o_4_7[4];
    data_i_4_8[4] = data_o_4_9[3];
    valid_i_4_8[4] = valid_o_4_9[3];
    ready_i_4_8[4] = ready_o_4_9[3];
    data_i_4_8[1] = data_o_3_8[2];
    valid_i_4_8[1] = valid_o_3_8[2];
    ready_i_4_8[1] = ready_o_3_8[2];
    data_i_4_8[2] = data_o_5_8[1];
    valid_i_4_8[2] = valid_o_5_8[1];
    ready_i_4_8[2] = ready_o_5_8[1];
    data_i_4_8[0] = data_i[4][8];
    valid_i_4_8[0] = valid_i[4][8];
    ready_i_4_8[0] = ready_i[4][8];
end


/*Router 4,9*/    
merge_router #(
    .input_mask                     (input_mask_4_9),
    .output_sel                     (output_sel_4_9)
)router94(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_4_9),
    .valid_i                        (valid_i_4_9),
    .ready_o                        (ready_o_4_9),
    .data_o                         (data_o_4_9),
    .valid_o                        (valid_o_4_9),
    .ready_i                        (ready_i_4_9)
);


always@(*) begin
    data_i_4_9[3] = data_o_4_8[4];
    valid_i_4_9[3] = valid_o_4_8[4];
    ready_i_4_9[3] = ready_o_4_8[4];
    data_i_4_9[4] = data_o_4_10[3];
    valid_i_4_9[4] = valid_o_4_10[3];
    ready_i_4_9[4] = ready_o_4_10[3];
    data_i_4_9[1] = data_o_3_9[2];
    valid_i_4_9[1] = valid_o_3_9[2];
    ready_i_4_9[1] = ready_o_3_9[2];
    data_i_4_9[2] = data_o_5_9[1];
    valid_i_4_9[2] = valid_o_5_9[1];
    ready_i_4_9[2] = ready_o_5_9[1];
    data_i_4_9[0] = data_i[4][9];
    valid_i_4_9[0] = valid_i[4][9];
    ready_i_4_9[0] = ready_i[4][9];
end


/*Router 4,10*/    
merge_router #(
    .input_mask                     (input_mask_4_10),
    .output_sel                     (output_sel_4_10)
)router104(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_4_10),
    .valid_i                        (valid_i_4_10),
    .ready_o                        (ready_o_4_10),
    .data_o                         (data_o_4_10),
    .valid_o                        (valid_o_4_10),
    .ready_i                        (ready_i_4_10)
);


always@(*) begin
    data_i_4_10[3] = data_o_4_9[4];
    valid_i_4_10[3] = valid_o_4_9[4];
    ready_i_4_10[3] = ready_o_4_9[4];
    data_i_4_10[4] = data_o_4_11[3];
    valid_i_4_10[4] = valid_o_4_11[3];
    ready_i_4_10[4] = ready_o_4_11[3];
    data_i_4_10[1] = data_o_3_10[2];
    valid_i_4_10[1] = valid_o_3_10[2];
    ready_i_4_10[1] = ready_o_3_10[2];
    data_i_4_10[2] = data_o_5_10[1];
    valid_i_4_10[2] = valid_o_5_10[1];
    ready_i_4_10[2] = ready_o_5_10[1];
    data_i_4_10[0] = data_i[4][10];
    valid_i_4_10[0] = valid_i[4][10];
    ready_i_4_10[0] = ready_i[4][10];
end


/*Router 4,11*/    
merge_router #(
    .input_mask                     (input_mask_4_11),
    .output_sel                     (output_sel_4_11)
)router114(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_4_11),
    .valid_i                        (valid_i_4_11),
    .ready_o                        (ready_o_4_11),
    .data_o                         (data_o_4_11),
    .valid_o                        (valid_o_4_11),
    .ready_i                        (ready_i_4_11)
);


always@(*) begin
    data_i_4_11[3] = data_o_4_10[4];
    valid_i_4_11[3] = valid_o_4_10[4];
    ready_i_4_11[3] = ready_o_4_10[4];
    data_i_4_11[4] = data_o_4_12[3];
    valid_i_4_11[4] = valid_o_4_12[3];
    ready_i_4_11[4] = ready_o_4_12[3];
    data_i_4_11[1] = data_o_3_11[2];
    valid_i_4_11[1] = valid_o_3_11[2];
    ready_i_4_11[1] = ready_o_3_11[2];
    data_i_4_11[2] = data_o_5_11[1];
    valid_i_4_11[2] = valid_o_5_11[1];
    ready_i_4_11[2] = ready_o_5_11[1];
    data_i_4_11[0] = data_i[4][11];
    valid_i_4_11[0] = valid_i[4][11];
    ready_i_4_11[0] = ready_i[4][11];
end


/*Router 4,12*/    
merge_router #(
    .input_mask                     (input_mask_4_12),
    .output_sel                     (output_sel_4_12)
)router124(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_4_12),
    .valid_i                        (valid_i_4_12),
    .ready_o                        (ready_o_4_12),
    .data_o                         (data_o_4_12),
    .valid_o                        (valid_o_4_12),
    .ready_i                        (ready_i_4_12)
);


always@(*) begin
    data_i_4_12[3] = data_o_4_11[4];
    valid_i_4_12[3] = valid_o_4_11[4];
    ready_i_4_12[3] = ready_o_4_11[4];
    data_i_4_12[4] = data_o_4_13[3];
    valid_i_4_12[4] = valid_o_4_13[3];
    ready_i_4_12[4] = ready_o_4_13[3];
    data_i_4_12[1] = data_o_3_12[2];
    valid_i_4_12[1] = valid_o_3_12[2];
    ready_i_4_12[1] = ready_o_3_12[2];
    data_i_4_12[2] = data_o_5_12[1];
    valid_i_4_12[2] = valid_o_5_12[1];
    ready_i_4_12[2] = ready_o_5_12[1];
    data_i_4_12[0] = data_i[4][12];
    valid_i_4_12[0] = valid_i[4][12];
    ready_i_4_12[0] = ready_i[4][12];
end


/*Router 4,13*/    
merge_router #(
    .input_mask                     (input_mask_4_13),
    .output_sel                     (output_sel_4_13)
)router134(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_4_13),
    .valid_i                        (valid_i_4_13),
    .ready_o                        (ready_o_4_13),
    .data_o                         (data_o_4_13),
    .valid_o                        (valid_o_4_13),
    .ready_i                        (ready_i_4_13)
);


always@(*) begin
    data_i_4_13[3] = data_o_4_12[4];
    valid_i_4_13[3] = valid_o_4_12[4];
    ready_i_4_13[3] = ready_o_4_12[4];
    data_i_4_13[4] = data_o_4_14[3];
    valid_i_4_13[4] = valid_o_4_14[3];
    ready_i_4_13[4] = ready_o_4_14[3];
    data_i_4_13[1] = data_o_3_13[2];
    valid_i_4_13[1] = valid_o_3_13[2];
    ready_i_4_13[1] = ready_o_3_13[2];
    data_i_4_13[2] = data_o_5_13[1];
    valid_i_4_13[2] = valid_o_5_13[1];
    ready_i_4_13[2] = ready_o_5_13[1];
    data_i_4_13[0] = data_i[4][13];
    valid_i_4_13[0] = valid_i[4][13];
    ready_i_4_13[0] = ready_i[4][13];
end


/*Router 4,14*/    
merge_router #(
    .input_mask                     (input_mask_4_14),
    .output_sel                     (output_sel_4_14)
)router144(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_4_14),
    .valid_i                        (valid_i_4_14),
    .ready_o                        (ready_o_4_14),
    .data_o                         (data_o_4_14),
    .valid_o                        (valid_o_4_14),
    .ready_i                        (ready_i_4_14)
);


always@(*) begin
    data_i_4_14[3] = data_o_4_13[4];
    valid_i_4_14[3] = valid_o_4_13[4];
    ready_i_4_14[3] = ready_o_4_13[4];
    data_i_4_14[4] = data_o_4_15[3];
    valid_i_4_14[4] = valid_o_4_15[3];
    ready_i_4_14[4] = ready_o_4_15[3];
    data_i_4_14[1] = data_o_3_14[2];
    valid_i_4_14[1] = valid_o_3_14[2];
    ready_i_4_14[1] = ready_o_3_14[2];
    data_i_4_14[2] = data_o_5_14[1];
    valid_i_4_14[2] = valid_o_5_14[1];
    ready_i_4_14[2] = ready_o_5_14[1];
    data_i_4_14[0] = data_i[4][14];
    valid_i_4_14[0] = valid_i[4][14];
    ready_i_4_14[0] = ready_i[4][14];
end


/*Router 4,15*/    
merge_router #(
    .input_mask                     (input_mask_4_15),
    .output_sel                     (output_sel_4_15)
)router154(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_4_15),
    .valid_i                        (valid_i_4_15),
    .ready_o                        (ready_o_4_15),
    .data_o                         (data_o_4_15),
    .valid_o                        (valid_o_4_15),
    .ready_i                        (ready_i_4_15)
);


always@(*) begin
    data_i_4_15[3] = data_o_4_14[4];
    valid_i_4_15[3] = valid_o_4_14[4];
    ready_i_4_15[3] = ready_o_4_14[4];
    data_i_4_15[4] = data_o_4_16[3];
    valid_i_4_15[4] = valid_o_4_16[3];
    ready_i_4_15[4] = ready_o_4_16[3];
    data_i_4_15[1] = data_o_3_15[2];
    valid_i_4_15[1] = valid_o_3_15[2];
    ready_i_4_15[1] = ready_o_3_15[2];
    data_i_4_15[2] = data_o_5_15[1];
    valid_i_4_15[2] = valid_o_5_15[1];
    ready_i_4_15[2] = ready_o_5_15[1];
    data_i_4_15[0] = data_i[4][15];
    valid_i_4_15[0] = valid_i[4][15];
    ready_i_4_15[0] = ready_i[4][15];
end


/*Router 4,16*/    
merge_router #(
    .input_mask                     (input_mask_4_16),
    .output_sel                     (output_sel_4_16)
)router164(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_4_16),
    .valid_i                        (valid_i_4_16),
    .ready_o                        (ready_o_4_16),
    .data_o                         (data_o_4_16),
    .valid_o                        (valid_o_4_16),
    .ready_i                        (ready_i_4_16)
);


always@(*) begin
    data_i_4_16[3] = data_o_4_15[4];
    valid_i_4_16[3] = valid_o_4_15[4];
    ready_i_4_16[3] = ready_o_4_15[4];
    data_i_4_16[4] = data_o_4_17[3];
    valid_i_4_16[4] = valid_o_4_17[3];
    ready_i_4_16[4] = ready_o_4_17[3];
    data_i_4_16[1] = data_o_3_16[2];
    valid_i_4_16[1] = valid_o_3_16[2];
    ready_i_4_16[1] = ready_o_3_16[2];
    data_i_4_16[2] = data_o_5_16[1];
    valid_i_4_16[2] = valid_o_5_16[1];
    ready_i_4_16[2] = ready_o_5_16[1];
    data_i_4_16[0] = data_i[4][16];
    valid_i_4_16[0] = valid_i[4][16];
    ready_i_4_16[0] = ready_i[4][16];
end


/*Router 4,17*/    
merge_router #(
    .input_mask                     (input_mask_4_17),
    .output_sel                     (output_sel_4_17)
)router174(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_4_17),
    .valid_i                        (valid_i_4_17),
    .ready_o                        (ready_o_4_17),
    .data_o                         (data_o_4_17),
    .valid_o                        (valid_o_4_17),
    .ready_i                        (ready_i_4_17)
);


always@(*) begin
    data_i_4_17[3] = data_o_4_16[4];
    valid_i_4_17[3] = valid_o_4_16[4];
    ready_i_4_17[3] = ready_o_4_16[4];
    data_i_4_17[4] = data_o_4_18[3];
    valid_i_4_17[4] = valid_o_4_18[3];
    ready_i_4_17[4] = ready_o_4_18[3];
    data_i_4_17[1] = data_o_3_17[2];
    valid_i_4_17[1] = valid_o_3_17[2];
    ready_i_4_17[1] = ready_o_3_17[2];
    data_i_4_17[2] = data_o_5_17[1];
    valid_i_4_17[2] = valid_o_5_17[1];
    ready_i_4_17[2] = ready_o_5_17[1];
    data_i_4_17[0] = data_i[4][17];
    valid_i_4_17[0] = valid_i[4][17];
    ready_i_4_17[0] = ready_i[4][17];
end


/*Router 4,18*/    
merge_router #(
    .input_mask                     (input_mask_4_18),
    .output_sel                     (output_sel_4_18)
)router184(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_4_18),
    .valid_i                        (valid_i_4_18),
    .ready_o                        (ready_o_4_18),
    .data_o                         (data_o_4_18),
    .valid_o                        (valid_o_4_18),
    .ready_i                        (ready_i_4_18)
);


always@(*) begin
    data_i_4_18[3] = data_o_4_17[4];
    valid_i_4_18[3] = valid_o_4_17[4];
    ready_i_4_18[3] = ready_o_4_17[4];
    data_i_4_18[4] = data_o_4_19[3];
    valid_i_4_18[4] = valid_o_4_19[3];
    ready_i_4_18[4] = ready_o_4_19[3];
    data_i_4_18[1] = data_o_3_18[2];
    valid_i_4_18[1] = valid_o_3_18[2];
    ready_i_4_18[1] = ready_o_3_18[2];
    data_i_4_18[2] = data_o_5_18[1];
    valid_i_4_18[2] = valid_o_5_18[1];
    ready_i_4_18[2] = ready_o_5_18[1];
    data_i_4_18[0] = data_i[4][18];
    valid_i_4_18[0] = valid_i[4][18];
    ready_i_4_18[0] = ready_i[4][18];
end


/*Router 4,19*/    
merge_router #(
    .input_mask                     (input_mask_4_19),
    .output_sel                     (output_sel_4_19)
)router194(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_4_19),
    .valid_i                        (valid_i_4_19),
    .ready_o                        (ready_o_4_19),
    .data_o                         (data_o_4_19),
    .valid_o                        (valid_o_4_19),
    .ready_i                        (ready_i_4_19)
);


always@(*) begin
    data_i_4_19[3] = data_o_4_18[4];
    valid_i_4_19[3] = valid_o_4_18[4];
    ready_i_4_19[3] = ready_o_4_18[4];
    data_i_4_19[4] = data_o_4_20[3];
    valid_i_4_19[4] = valid_o_4_20[3];
    ready_i_4_19[4] = ready_o_4_20[3];
    data_i_4_19[1] = data_o_3_19[2];
    valid_i_4_19[1] = valid_o_3_19[2];
    ready_i_4_19[1] = ready_o_3_19[2];
    data_i_4_19[2] = data_o_5_19[1];
    valid_i_4_19[2] = valid_o_5_19[1];
    ready_i_4_19[2] = ready_o_5_19[1];
    data_i_4_19[0] = data_i[4][19];
    valid_i_4_19[0] = valid_i[4][19];
    ready_i_4_19[0] = ready_i[4][19];
end


/*Router 4,20*/    
merge_router #(
    .input_mask                     (input_mask_4_20),
    .output_sel                     (output_sel_4_20)
)router204(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_4_20),
    .valid_i                        (valid_i_4_20),
    .ready_o                        (ready_o_4_20),
    .data_o                         (data_o_4_20),
    .valid_o                        (valid_o_4_20),
    .ready_i                        (ready_i_4_20)
);


always@(*) begin
    data_i_4_20[3] = data_o_4_19[4];
    valid_i_4_20[3] = valid_o_4_19[4];
    ready_i_4_20[3] = ready_o_4_19[4];
    data_i_4_20[4] = data_o_4_21[3];
    valid_i_4_20[4] = valid_o_4_21[3];
    ready_i_4_20[4] = ready_o_4_21[3];
    data_i_4_20[1] = data_o_3_20[2];
    valid_i_4_20[1] = valid_o_3_20[2];
    ready_i_4_20[1] = ready_o_3_20[2];
    data_i_4_20[2] = data_o_5_20[1];
    valid_i_4_20[2] = valid_o_5_20[1];
    ready_i_4_20[2] = ready_o_5_20[1];
    data_i_4_20[0] = data_i[4][20];
    valid_i_4_20[0] = valid_i[4][20];
    ready_i_4_20[0] = ready_i[4][20];
end


/*Router 4,21*/    
merge_router #(
    .input_mask                     (input_mask_4_21),
    .output_sel                     (output_sel_4_21)
)router214(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_4_21),
    .valid_i                        (valid_i_4_21),
    .ready_o                        (ready_o_4_21),
    .data_o                         (data_o_4_21),
    .valid_o                        (valid_o_4_21),
    .ready_i                        (ready_i_4_21)
);


always@(*) begin
    data_i_4_21[3] = data_o_4_20[4];
    valid_i_4_21[3] = valid_o_4_20[4];
    ready_i_4_21[3] = ready_o_4_20[4];
    data_i_4_21[4] = data_o_4_22[3];
    valid_i_4_21[4] = valid_o_4_22[3];
    ready_i_4_21[4] = ready_o_4_22[3];
    data_i_4_21[1] = data_o_3_21[2];
    valid_i_4_21[1] = valid_o_3_21[2];
    ready_i_4_21[1] = ready_o_3_21[2];
    data_i_4_21[2] = data_o_5_21[1];
    valid_i_4_21[2] = valid_o_5_21[1];
    ready_i_4_21[2] = ready_o_5_21[1];
    data_i_4_21[0] = data_i[4][21];
    valid_i_4_21[0] = valid_i[4][21];
    ready_i_4_21[0] = ready_i[4][21];
end


/*Router 4,22*/    
merge_router #(
    .input_mask                     (input_mask_4_22),
    .output_sel                     (output_sel_4_22)
)router224(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_4_22),
    .valid_i                        (valid_i_4_22),
    .ready_o                        (ready_o_4_22),
    .data_o                         (data_o_4_22),
    .valid_o                        (valid_o_4_22),
    .ready_i                        (ready_i_4_22)
);


always@(*) begin
    data_i_4_22[3] = data_o_4_21[4];
    valid_i_4_22[3] = valid_o_4_21[4];
    ready_i_4_22[3] = ready_o_4_21[4];
    data_i_4_22[4] = data_o_4_23[3];
    valid_i_4_22[4] = valid_o_4_23[3];
    ready_i_4_22[4] = ready_o_4_23[3];
    data_i_4_22[1] = data_o_3_22[2];
    valid_i_4_22[1] = valid_o_3_22[2];
    ready_i_4_22[1] = ready_o_3_22[2];
    data_i_4_22[2] = data_o_5_22[1];
    valid_i_4_22[2] = valid_o_5_22[1];
    ready_i_4_22[2] = ready_o_5_22[1];
    data_i_4_22[0] = data_i[4][22];
    valid_i_4_22[0] = valid_i[4][22];
    ready_i_4_22[0] = ready_i[4][22];
end


/*Router 4,23*/    
merge_router #(
    .input_mask                     (input_mask_4_23),
    .output_sel                     (output_sel_4_23)
)router234(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_4_23),
    .valid_i                        (valid_i_4_23),
    .ready_o                        (ready_o_4_23),
    .data_o                         (data_o_4_23),
    .valid_o                        (valid_o_4_23),
    .ready_i                        (ready_i_4_23)
);


always@(*) begin
    data_i_4_23[3] = data_o_4_22[4];
    valid_i_4_23[3] = valid_o_4_22[4];
    ready_i_4_23[3] = ready_o_4_22[4];
    data_i_4_23[4] = data_o_4_24[3];
    valid_i_4_23[4] = valid_o_4_24[3];
    ready_i_4_23[4] = ready_o_4_24[3];
    data_i_4_23[1] = data_o_3_23[2];
    valid_i_4_23[1] = valid_o_3_23[2];
    ready_i_4_23[1] = ready_o_3_23[2];
    data_i_4_23[2] = data_o_5_23[1];
    valid_i_4_23[2] = valid_o_5_23[1];
    ready_i_4_23[2] = ready_o_5_23[1];
    data_i_4_23[0] = data_i[4][23];
    valid_i_4_23[0] = valid_i[4][23];
    ready_i_4_23[0] = ready_i[4][23];
end


/*Router 4,24*/    
merge_router #(
    .input_mask                     (input_mask_4_24),
    .output_sel                     (output_sel_4_24)
)router244(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_4_24),
    .valid_i                        (valid_i_4_24),
    .ready_o                        (ready_o_4_24),
    .data_o                         (data_o_4_24),
    .valid_o                        (valid_o_4_24),
    .ready_i                        (ready_i_4_24)
);


always@(*) begin
    data_i_4_24[3] = data_o_4_23[4];
    valid_i_4_24[3] = valid_o_4_23[4];
    ready_i_4_24[3] = ready_o_4_23[4];
    data_i_4_24[1] = data_o_3_24[2];
    valid_i_4_24[1] = valid_o_3_24[2];
    ready_i_4_24[1] = ready_o_3_24[2];
    data_i_4_24[2] = data_o_5_24[1];
    valid_i_4_24[2] = valid_o_5_24[1];
    ready_i_4_24[2] = ready_o_5_24[1];
    data_i_4_24[0] = data_i[4][24];
    valid_i_4_24[0] = valid_i[4][24];
    ready_i_4_24[0] = ready_i[4][24];
end


/*Router 5,0*/    
merge_router #(
    .input_mask                     (input_mask_5_0),
    .output_sel                     (output_sel_5_0)
)router5(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_5_0),
    .valid_i                        (valid_i_5_0),
    .ready_o                        (ready_o_5_0),
    .data_o                         (data_o_5_0),
    .valid_o                        (valid_o_5_0),
    .ready_i                        (ready_i_5_0)
);


always@(*) begin
    data_i_5_0[4] = data_o_5_1[3];
    valid_i_5_0[4] = valid_o_5_1[3];
    ready_i_5_0[4] = ready_o_5_1[3];
    data_i_5_0[1] = data_o_4_0[2];
    valid_i_5_0[1] = valid_o_4_0[2];
    ready_i_5_0[1] = ready_o_4_0[2];
    data_i_5_0[2] = data_o_6_0[1];
    valid_i_5_0[2] = valid_o_6_0[1];
    ready_i_5_0[2] = ready_o_6_0[1];
    data_i_5_0[0] = data_i[5][0];
    valid_i_5_0[0] = valid_i[5][0];
    ready_i_5_0[0] = ready_i[5][0];
end


/*Router 5,1*/    
merge_router #(
    .input_mask                     (input_mask_5_1),
    .output_sel                     (output_sel_5_1)
)router15(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_5_1),
    .valid_i                        (valid_i_5_1),
    .ready_o                        (ready_o_5_1),
    .data_o                         (data_o_5_1),
    .valid_o                        (valid_o_5_1),
    .ready_i                        (ready_i_5_1)
);


always@(*) begin
    data_i_5_1[3] = data_o_5_0[4];
    valid_i_5_1[3] = valid_o_5_0[4];
    ready_i_5_1[3] = ready_o_5_0[4];
    data_i_5_1[4] = data_o_5_2[3];
    valid_i_5_1[4] = valid_o_5_2[3];
    ready_i_5_1[4] = ready_o_5_2[3];
    data_i_5_1[1] = data_o_4_1[2];
    valid_i_5_1[1] = valid_o_4_1[2];
    ready_i_5_1[1] = ready_o_4_1[2];
    data_i_5_1[2] = data_o_6_1[1];
    valid_i_5_1[2] = valid_o_6_1[1];
    ready_i_5_1[2] = ready_o_6_1[1];
    data_i_5_1[0] = data_i[5][1];
    valid_i_5_1[0] = valid_i[5][1];
    ready_i_5_1[0] = ready_i[5][1];
end


/*Router 5,2*/    
merge_router #(
    .input_mask                     (input_mask_5_2),
    .output_sel                     (output_sel_5_2)
)router25(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_5_2),
    .valid_i                        (valid_i_5_2),
    .ready_o                        (ready_o_5_2),
    .data_o                         (data_o_5_2),
    .valid_o                        (valid_o_5_2),
    .ready_i                        (ready_i_5_2)
);


always@(*) begin
    data_i_5_2[3] = data_o_5_1[4];
    valid_i_5_2[3] = valid_o_5_1[4];
    ready_i_5_2[3] = ready_o_5_1[4];
    data_i_5_2[4] = data_o_5_3[3];
    valid_i_5_2[4] = valid_o_5_3[3];
    ready_i_5_2[4] = ready_o_5_3[3];
    data_i_5_2[1] = data_o_4_2[2];
    valid_i_5_2[1] = valid_o_4_2[2];
    ready_i_5_2[1] = ready_o_4_2[2];
    data_i_5_2[2] = data_o_6_2[1];
    valid_i_5_2[2] = valid_o_6_2[1];
    ready_i_5_2[2] = ready_o_6_2[1];
    data_i_5_2[0] = data_i[5][2];
    valid_i_5_2[0] = valid_i[5][2];
    ready_i_5_2[0] = ready_i[5][2];
end


/*Router 5,3*/    
merge_router #(
    .input_mask                     (input_mask_5_3),
    .output_sel                     (output_sel_5_3)
)router35(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_5_3),
    .valid_i                        (valid_i_5_3),
    .ready_o                        (ready_o_5_3),
    .data_o                         (data_o_5_3),
    .valid_o                        (valid_o_5_3),
    .ready_i                        (ready_i_5_3)
);


always@(*) begin
    data_i_5_3[3] = data_o_5_2[4];
    valid_i_5_3[3] = valid_o_5_2[4];
    ready_i_5_3[3] = ready_o_5_2[4];
    data_i_5_3[4] = data_o_5_4[3];
    valid_i_5_3[4] = valid_o_5_4[3];
    ready_i_5_3[4] = ready_o_5_4[3];
    data_i_5_3[1] = data_o_4_3[2];
    valid_i_5_3[1] = valid_o_4_3[2];
    ready_i_5_3[1] = ready_o_4_3[2];
    data_i_5_3[2] = data_o_6_3[1];
    valid_i_5_3[2] = valid_o_6_3[1];
    ready_i_5_3[2] = ready_o_6_3[1];
    data_i_5_3[0] = data_i[5][3];
    valid_i_5_3[0] = valid_i[5][3];
    ready_i_5_3[0] = ready_i[5][3];
end


/*Router 5,4*/    
merge_router #(
    .input_mask                     (input_mask_5_4),
    .output_sel                     (output_sel_5_4)
)router45(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_5_4),
    .valid_i                        (valid_i_5_4),
    .ready_o                        (ready_o_5_4),
    .data_o                         (data_o_5_4),
    .valid_o                        (valid_o_5_4),
    .ready_i                        (ready_i_5_4)
);


always@(*) begin
    data_i_5_4[3] = data_o_5_3[4];
    valid_i_5_4[3] = valid_o_5_3[4];
    ready_i_5_4[3] = ready_o_5_3[4];
    data_i_5_4[4] = data_o_5_5[3];
    valid_i_5_4[4] = valid_o_5_5[3];
    ready_i_5_4[4] = ready_o_5_5[3];
    data_i_5_4[1] = data_o_4_4[2];
    valid_i_5_4[1] = valid_o_4_4[2];
    ready_i_5_4[1] = ready_o_4_4[2];
    data_i_5_4[2] = data_o_6_4[1];
    valid_i_5_4[2] = valid_o_6_4[1];
    ready_i_5_4[2] = ready_o_6_4[1];
    data_i_5_4[0] = data_i[5][4];
    valid_i_5_4[0] = valid_i[5][4];
    ready_i_5_4[0] = ready_i[5][4];
end


/*Router 5,5*/    
merge_router #(
    .input_mask                     (input_mask_5_5),
    .output_sel                     (output_sel_5_5)
)router55(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_5_5),
    .valid_i                        (valid_i_5_5),
    .ready_o                        (ready_o_5_5),
    .data_o                         (data_o_5_5),
    .valid_o                        (valid_o_5_5),
    .ready_i                        (ready_i_5_5)
);


always@(*) begin
    data_i_5_5[3] = data_o_5_4[4];
    valid_i_5_5[3] = valid_o_5_4[4];
    ready_i_5_5[3] = ready_o_5_4[4];
    data_i_5_5[4] = data_o_5_6[3];
    valid_i_5_5[4] = valid_o_5_6[3];
    ready_i_5_5[4] = ready_o_5_6[3];
    data_i_5_5[1] = data_o_4_5[2];
    valid_i_5_5[1] = valid_o_4_5[2];
    ready_i_5_5[1] = ready_o_4_5[2];
    data_i_5_5[2] = data_o_6_5[1];
    valid_i_5_5[2] = valid_o_6_5[1];
    ready_i_5_5[2] = ready_o_6_5[1];
    data_i_5_5[0] = data_i[5][5];
    valid_i_5_5[0] = valid_i[5][5];
    ready_i_5_5[0] = ready_i[5][5];
end


/*Router 5,6*/    
merge_router #(
    .input_mask                     (input_mask_5_6),
    .output_sel                     (output_sel_5_6)
)router65(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_5_6),
    .valid_i                        (valid_i_5_6),
    .ready_o                        (ready_o_5_6),
    .data_o                         (data_o_5_6),
    .valid_o                        (valid_o_5_6),
    .ready_i                        (ready_i_5_6)
);


always@(*) begin
    data_i_5_6[3] = data_o_5_5[4];
    valid_i_5_6[3] = valid_o_5_5[4];
    ready_i_5_6[3] = ready_o_5_5[4];
    data_i_5_6[4] = data_o_5_7[3];
    valid_i_5_6[4] = valid_o_5_7[3];
    ready_i_5_6[4] = ready_o_5_7[3];
    data_i_5_6[1] = data_o_4_6[2];
    valid_i_5_6[1] = valid_o_4_6[2];
    ready_i_5_6[1] = ready_o_4_6[2];
    data_i_5_6[2] = data_o_6_6[1];
    valid_i_5_6[2] = valid_o_6_6[1];
    ready_i_5_6[2] = ready_o_6_6[1];
    data_i_5_6[0] = data_i[5][6];
    valid_i_5_6[0] = valid_i[5][6];
    ready_i_5_6[0] = ready_i[5][6];
end


/*Router 5,7*/    
merge_router #(
    .input_mask                     (input_mask_5_7),
    .output_sel                     (output_sel_5_7)
)router75(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_5_7),
    .valid_i                        (valid_i_5_7),
    .ready_o                        (ready_o_5_7),
    .data_o                         (data_o_5_7),
    .valid_o                        (valid_o_5_7),
    .ready_i                        (ready_i_5_7)
);


always@(*) begin
    data_i_5_7[3] = data_o_5_6[4];
    valid_i_5_7[3] = valid_o_5_6[4];
    ready_i_5_7[3] = ready_o_5_6[4];
    data_i_5_7[4] = data_o_5_8[3];
    valid_i_5_7[4] = valid_o_5_8[3];
    ready_i_5_7[4] = ready_o_5_8[3];
    data_i_5_7[1] = data_o_4_7[2];
    valid_i_5_7[1] = valid_o_4_7[2];
    ready_i_5_7[1] = ready_o_4_7[2];
    data_i_5_7[2] = data_o_6_7[1];
    valid_i_5_7[2] = valid_o_6_7[1];
    ready_i_5_7[2] = ready_o_6_7[1];
    data_i_5_7[0] = data_i[5][7];
    valid_i_5_7[0] = valid_i[5][7];
    ready_i_5_7[0] = ready_i[5][7];
end


/*Router 5,8*/    
merge_router #(
    .input_mask                     (input_mask_5_8),
    .output_sel                     (output_sel_5_8)
)router85(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_5_8),
    .valid_i                        (valid_i_5_8),
    .ready_o                        (ready_o_5_8),
    .data_o                         (data_o_5_8),
    .valid_o                        (valid_o_5_8),
    .ready_i                        (ready_i_5_8)
);


always@(*) begin
    data_i_5_8[3] = data_o_5_7[4];
    valid_i_5_8[3] = valid_o_5_7[4];
    ready_i_5_8[3] = ready_o_5_7[4];
    data_i_5_8[4] = data_o_5_9[3];
    valid_i_5_8[4] = valid_o_5_9[3];
    ready_i_5_8[4] = ready_o_5_9[3];
    data_i_5_8[1] = data_o_4_8[2];
    valid_i_5_8[1] = valid_o_4_8[2];
    ready_i_5_8[1] = ready_o_4_8[2];
    data_i_5_8[2] = data_o_6_8[1];
    valid_i_5_8[2] = valid_o_6_8[1];
    ready_i_5_8[2] = ready_o_6_8[1];
    data_i_5_8[0] = data_i[5][8];
    valid_i_5_8[0] = valid_i[5][8];
    ready_i_5_8[0] = ready_i[5][8];
end


/*Router 5,9*/    
merge_router #(
    .input_mask                     (input_mask_5_9),
    .output_sel                     (output_sel_5_9)
)router95(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_5_9),
    .valid_i                        (valid_i_5_9),
    .ready_o                        (ready_o_5_9),
    .data_o                         (data_o_5_9),
    .valid_o                        (valid_o_5_9),
    .ready_i                        (ready_i_5_9)
);


always@(*) begin
    data_i_5_9[3] = data_o_5_8[4];
    valid_i_5_9[3] = valid_o_5_8[4];
    ready_i_5_9[3] = ready_o_5_8[4];
    data_i_5_9[4] = data_o_5_10[3];
    valid_i_5_9[4] = valid_o_5_10[3];
    ready_i_5_9[4] = ready_o_5_10[3];
    data_i_5_9[1] = data_o_4_9[2];
    valid_i_5_9[1] = valid_o_4_9[2];
    ready_i_5_9[1] = ready_o_4_9[2];
    data_i_5_9[2] = data_o_6_9[1];
    valid_i_5_9[2] = valid_o_6_9[1];
    ready_i_5_9[2] = ready_o_6_9[1];
    data_i_5_9[0] = data_i[5][9];
    valid_i_5_9[0] = valid_i[5][9];
    ready_i_5_9[0] = ready_i[5][9];
end


/*Router 5,10*/    
merge_router #(
    .input_mask                     (input_mask_5_10),
    .output_sel                     (output_sel_5_10)
)router105(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_5_10),
    .valid_i                        (valid_i_5_10),
    .ready_o                        (ready_o_5_10),
    .data_o                         (data_o_5_10),
    .valid_o                        (valid_o_5_10),
    .ready_i                        (ready_i_5_10)
);


always@(*) begin
    data_i_5_10[3] = data_o_5_9[4];
    valid_i_5_10[3] = valid_o_5_9[4];
    ready_i_5_10[3] = ready_o_5_9[4];
    data_i_5_10[4] = data_o_5_11[3];
    valid_i_5_10[4] = valid_o_5_11[3];
    ready_i_5_10[4] = ready_o_5_11[3];
    data_i_5_10[1] = data_o_4_10[2];
    valid_i_5_10[1] = valid_o_4_10[2];
    ready_i_5_10[1] = ready_o_4_10[2];
    data_i_5_10[2] = data_o_6_10[1];
    valid_i_5_10[2] = valid_o_6_10[1];
    ready_i_5_10[2] = ready_o_6_10[1];
    data_i_5_10[0] = data_i[5][10];
    valid_i_5_10[0] = valid_i[5][10];
    ready_i_5_10[0] = ready_i[5][10];
end


/*Router 5,11*/    
merge_router #(
    .input_mask                     (input_mask_5_11),
    .output_sel                     (output_sel_5_11)
)router115(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_5_11),
    .valid_i                        (valid_i_5_11),
    .ready_o                        (ready_o_5_11),
    .data_o                         (data_o_5_11),
    .valid_o                        (valid_o_5_11),
    .ready_i                        (ready_i_5_11)
);


always@(*) begin
    data_i_5_11[3] = data_o_5_10[4];
    valid_i_5_11[3] = valid_o_5_10[4];
    ready_i_5_11[3] = ready_o_5_10[4];
    data_i_5_11[4] = data_o_5_12[3];
    valid_i_5_11[4] = valid_o_5_12[3];
    ready_i_5_11[4] = ready_o_5_12[3];
    data_i_5_11[1] = data_o_4_11[2];
    valid_i_5_11[1] = valid_o_4_11[2];
    ready_i_5_11[1] = ready_o_4_11[2];
    data_i_5_11[2] = data_o_6_11[1];
    valid_i_5_11[2] = valid_o_6_11[1];
    ready_i_5_11[2] = ready_o_6_11[1];
    data_i_5_11[0] = data_i[5][11];
    valid_i_5_11[0] = valid_i[5][11];
    ready_i_5_11[0] = ready_i[5][11];
end


/*Router 5,12*/    
merge_router #(
    .input_mask                     (input_mask_5_12),
    .output_sel                     (output_sel_5_12)
)router125(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_5_12),
    .valid_i                        (valid_i_5_12),
    .ready_o                        (ready_o_5_12),
    .data_o                         (data_o_5_12),
    .valid_o                        (valid_o_5_12),
    .ready_i                        (ready_i_5_12)
);


always@(*) begin
    data_i_5_12[3] = data_o_5_11[4];
    valid_i_5_12[3] = valid_o_5_11[4];
    ready_i_5_12[3] = ready_o_5_11[4];
    data_i_5_12[4] = data_o_5_13[3];
    valid_i_5_12[4] = valid_o_5_13[3];
    ready_i_5_12[4] = ready_o_5_13[3];
    data_i_5_12[1] = data_o_4_12[2];
    valid_i_5_12[1] = valid_o_4_12[2];
    ready_i_5_12[1] = ready_o_4_12[2];
    data_i_5_12[2] = data_o_6_12[1];
    valid_i_5_12[2] = valid_o_6_12[1];
    ready_i_5_12[2] = ready_o_6_12[1];
    data_i_5_12[0] = data_i[5][12];
    valid_i_5_12[0] = valid_i[5][12];
    ready_i_5_12[0] = ready_i[5][12];
end


/*Router 5,13*/    
merge_router #(
    .input_mask                     (input_mask_5_13),
    .output_sel                     (output_sel_5_13)
)router135(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_5_13),
    .valid_i                        (valid_i_5_13),
    .ready_o                        (ready_o_5_13),
    .data_o                         (data_o_5_13),
    .valid_o                        (valid_o_5_13),
    .ready_i                        (ready_i_5_13)
);


always@(*) begin
    data_i_5_13[3] = data_o_5_12[4];
    valid_i_5_13[3] = valid_o_5_12[4];
    ready_i_5_13[3] = ready_o_5_12[4];
    data_i_5_13[4] = data_o_5_14[3];
    valid_i_5_13[4] = valid_o_5_14[3];
    ready_i_5_13[4] = ready_o_5_14[3];
    data_i_5_13[1] = data_o_4_13[2];
    valid_i_5_13[1] = valid_o_4_13[2];
    ready_i_5_13[1] = ready_o_4_13[2];
    data_i_5_13[2] = data_o_6_13[1];
    valid_i_5_13[2] = valid_o_6_13[1];
    ready_i_5_13[2] = ready_o_6_13[1];
    data_i_5_13[0] = data_i[5][13];
    valid_i_5_13[0] = valid_i[5][13];
    ready_i_5_13[0] = ready_i[5][13];
end


/*Router 5,14*/    
merge_router #(
    .input_mask                     (input_mask_5_14),
    .output_sel                     (output_sel_5_14)
)router145(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_5_14),
    .valid_i                        (valid_i_5_14),
    .ready_o                        (ready_o_5_14),
    .data_o                         (data_o_5_14),
    .valid_o                        (valid_o_5_14),
    .ready_i                        (ready_i_5_14)
);


always@(*) begin
    data_i_5_14[3] = data_o_5_13[4];
    valid_i_5_14[3] = valid_o_5_13[4];
    ready_i_5_14[3] = ready_o_5_13[4];
    data_i_5_14[4] = data_o_5_15[3];
    valid_i_5_14[4] = valid_o_5_15[3];
    ready_i_5_14[4] = ready_o_5_15[3];
    data_i_5_14[1] = data_o_4_14[2];
    valid_i_5_14[1] = valid_o_4_14[2];
    ready_i_5_14[1] = ready_o_4_14[2];
    data_i_5_14[2] = data_o_6_14[1];
    valid_i_5_14[2] = valid_o_6_14[1];
    ready_i_5_14[2] = ready_o_6_14[1];
    data_i_5_14[0] = data_i[5][14];
    valid_i_5_14[0] = valid_i[5][14];
    ready_i_5_14[0] = ready_i[5][14];
end


/*Router 5,15*/    
merge_router #(
    .input_mask                     (input_mask_5_15),
    .output_sel                     (output_sel_5_15)
)router155(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_5_15),
    .valid_i                        (valid_i_5_15),
    .ready_o                        (ready_o_5_15),
    .data_o                         (data_o_5_15),
    .valid_o                        (valid_o_5_15),
    .ready_i                        (ready_i_5_15)
);


always@(*) begin
    data_i_5_15[3] = data_o_5_14[4];
    valid_i_5_15[3] = valid_o_5_14[4];
    ready_i_5_15[3] = ready_o_5_14[4];
    data_i_5_15[4] = data_o_5_16[3];
    valid_i_5_15[4] = valid_o_5_16[3];
    ready_i_5_15[4] = ready_o_5_16[3];
    data_i_5_15[1] = data_o_4_15[2];
    valid_i_5_15[1] = valid_o_4_15[2];
    ready_i_5_15[1] = ready_o_4_15[2];
    data_i_5_15[2] = data_o_6_15[1];
    valid_i_5_15[2] = valid_o_6_15[1];
    ready_i_5_15[2] = ready_o_6_15[1];
    data_i_5_15[0] = data_i[5][15];
    valid_i_5_15[0] = valid_i[5][15];
    ready_i_5_15[0] = ready_i[5][15];
end


/*Router 5,16*/    
merge_router #(
    .input_mask                     (input_mask_5_16),
    .output_sel                     (output_sel_5_16)
)router165(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_5_16),
    .valid_i                        (valid_i_5_16),
    .ready_o                        (ready_o_5_16),
    .data_o                         (data_o_5_16),
    .valid_o                        (valid_o_5_16),
    .ready_i                        (ready_i_5_16)
);


always@(*) begin
    data_i_5_16[3] = data_o_5_15[4];
    valid_i_5_16[3] = valid_o_5_15[4];
    ready_i_5_16[3] = ready_o_5_15[4];
    data_i_5_16[4] = data_o_5_17[3];
    valid_i_5_16[4] = valid_o_5_17[3];
    ready_i_5_16[4] = ready_o_5_17[3];
    data_i_5_16[1] = data_o_4_16[2];
    valid_i_5_16[1] = valid_o_4_16[2];
    ready_i_5_16[1] = ready_o_4_16[2];
    data_i_5_16[2] = data_o_6_16[1];
    valid_i_5_16[2] = valid_o_6_16[1];
    ready_i_5_16[2] = ready_o_6_16[1];
    data_i_5_16[0] = data_i[5][16];
    valid_i_5_16[0] = valid_i[5][16];
    ready_i_5_16[0] = ready_i[5][16];
end


/*Router 5,17*/    
merge_router #(
    .input_mask                     (input_mask_5_17),
    .output_sel                     (output_sel_5_17)
)router175(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_5_17),
    .valid_i                        (valid_i_5_17),
    .ready_o                        (ready_o_5_17),
    .data_o                         (data_o_5_17),
    .valid_o                        (valid_o_5_17),
    .ready_i                        (ready_i_5_17)
);


always@(*) begin
    data_i_5_17[3] = data_o_5_16[4];
    valid_i_5_17[3] = valid_o_5_16[4];
    ready_i_5_17[3] = ready_o_5_16[4];
    data_i_5_17[4] = data_o_5_18[3];
    valid_i_5_17[4] = valid_o_5_18[3];
    ready_i_5_17[4] = ready_o_5_18[3];
    data_i_5_17[1] = data_o_4_17[2];
    valid_i_5_17[1] = valid_o_4_17[2];
    ready_i_5_17[1] = ready_o_4_17[2];
    data_i_5_17[2] = data_o_6_17[1];
    valid_i_5_17[2] = valid_o_6_17[1];
    ready_i_5_17[2] = ready_o_6_17[1];
    data_i_5_17[0] = data_i[5][17];
    valid_i_5_17[0] = valid_i[5][17];
    ready_i_5_17[0] = ready_i[5][17];
end


/*Router 5,18*/    
merge_router #(
    .input_mask                     (input_mask_5_18),
    .output_sel                     (output_sel_5_18)
)router185(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_5_18),
    .valid_i                        (valid_i_5_18),
    .ready_o                        (ready_o_5_18),
    .data_o                         (data_o_5_18),
    .valid_o                        (valid_o_5_18),
    .ready_i                        (ready_i_5_18)
);


always@(*) begin
    data_i_5_18[3] = data_o_5_17[4];
    valid_i_5_18[3] = valid_o_5_17[4];
    ready_i_5_18[3] = ready_o_5_17[4];
    data_i_5_18[4] = data_o_5_19[3];
    valid_i_5_18[4] = valid_o_5_19[3];
    ready_i_5_18[4] = ready_o_5_19[3];
    data_i_5_18[1] = data_o_4_18[2];
    valid_i_5_18[1] = valid_o_4_18[2];
    ready_i_5_18[1] = ready_o_4_18[2];
    data_i_5_18[2] = data_o_6_18[1];
    valid_i_5_18[2] = valid_o_6_18[1];
    ready_i_5_18[2] = ready_o_6_18[1];
    data_i_5_18[0] = data_i[5][18];
    valid_i_5_18[0] = valid_i[5][18];
    ready_i_5_18[0] = ready_i[5][18];
end


/*Router 5,19*/    
merge_router #(
    .input_mask                     (input_mask_5_19),
    .output_sel                     (output_sel_5_19)
)router195(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_5_19),
    .valid_i                        (valid_i_5_19),
    .ready_o                        (ready_o_5_19),
    .data_o                         (data_o_5_19),
    .valid_o                        (valid_o_5_19),
    .ready_i                        (ready_i_5_19)
);


always@(*) begin
    data_i_5_19[3] = data_o_5_18[4];
    valid_i_5_19[3] = valid_o_5_18[4];
    ready_i_5_19[3] = ready_o_5_18[4];
    data_i_5_19[4] = data_o_5_20[3];
    valid_i_5_19[4] = valid_o_5_20[3];
    ready_i_5_19[4] = ready_o_5_20[3];
    data_i_5_19[1] = data_o_4_19[2];
    valid_i_5_19[1] = valid_o_4_19[2];
    ready_i_5_19[1] = ready_o_4_19[2];
    data_i_5_19[2] = data_o_6_19[1];
    valid_i_5_19[2] = valid_o_6_19[1];
    ready_i_5_19[2] = ready_o_6_19[1];
    data_i_5_19[0] = data_i[5][19];
    valid_i_5_19[0] = valid_i[5][19];
    ready_i_5_19[0] = ready_i[5][19];
end


/*Router 5,20*/    
merge_router #(
    .input_mask                     (input_mask_5_20),
    .output_sel                     (output_sel_5_20)
)router205(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_5_20),
    .valid_i                        (valid_i_5_20),
    .ready_o                        (ready_o_5_20),
    .data_o                         (data_o_5_20),
    .valid_o                        (valid_o_5_20),
    .ready_i                        (ready_i_5_20)
);


always@(*) begin
    data_i_5_20[3] = data_o_5_19[4];
    valid_i_5_20[3] = valid_o_5_19[4];
    ready_i_5_20[3] = ready_o_5_19[4];
    data_i_5_20[4] = data_o_5_21[3];
    valid_i_5_20[4] = valid_o_5_21[3];
    ready_i_5_20[4] = ready_o_5_21[3];
    data_i_5_20[1] = data_o_4_20[2];
    valid_i_5_20[1] = valid_o_4_20[2];
    ready_i_5_20[1] = ready_o_4_20[2];
    data_i_5_20[2] = data_o_6_20[1];
    valid_i_5_20[2] = valid_o_6_20[1];
    ready_i_5_20[2] = ready_o_6_20[1];
    data_i_5_20[0] = data_i[5][20];
    valid_i_5_20[0] = valid_i[5][20];
    ready_i_5_20[0] = ready_i[5][20];
end


/*Router 5,21*/    
merge_router #(
    .input_mask                     (input_mask_5_21),
    .output_sel                     (output_sel_5_21)
)router215(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_5_21),
    .valid_i                        (valid_i_5_21),
    .ready_o                        (ready_o_5_21),
    .data_o                         (data_o_5_21),
    .valid_o                        (valid_o_5_21),
    .ready_i                        (ready_i_5_21)
);


always@(*) begin
    data_i_5_21[3] = data_o_5_20[4];
    valid_i_5_21[3] = valid_o_5_20[4];
    ready_i_5_21[3] = ready_o_5_20[4];
    data_i_5_21[4] = data_o_5_22[3];
    valid_i_5_21[4] = valid_o_5_22[3];
    ready_i_5_21[4] = ready_o_5_22[3];
    data_i_5_21[1] = data_o_4_21[2];
    valid_i_5_21[1] = valid_o_4_21[2];
    ready_i_5_21[1] = ready_o_4_21[2];
    data_i_5_21[2] = data_o_6_21[1];
    valid_i_5_21[2] = valid_o_6_21[1];
    ready_i_5_21[2] = ready_o_6_21[1];
    data_i_5_21[0] = data_i[5][21];
    valid_i_5_21[0] = valid_i[5][21];
    ready_i_5_21[0] = ready_i[5][21];
end


/*Router 5,22*/    
merge_router #(
    .input_mask                     (input_mask_5_22),
    .output_sel                     (output_sel_5_22)
)router225(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_5_22),
    .valid_i                        (valid_i_5_22),
    .ready_o                        (ready_o_5_22),
    .data_o                         (data_o_5_22),
    .valid_o                        (valid_o_5_22),
    .ready_i                        (ready_i_5_22)
);


always@(*) begin
    data_i_5_22[3] = data_o_5_21[4];
    valid_i_5_22[3] = valid_o_5_21[4];
    ready_i_5_22[3] = ready_o_5_21[4];
    data_i_5_22[4] = data_o_5_23[3];
    valid_i_5_22[4] = valid_o_5_23[3];
    ready_i_5_22[4] = ready_o_5_23[3];
    data_i_5_22[1] = data_o_4_22[2];
    valid_i_5_22[1] = valid_o_4_22[2];
    ready_i_5_22[1] = ready_o_4_22[2];
    data_i_5_22[2] = data_o_6_22[1];
    valid_i_5_22[2] = valid_o_6_22[1];
    ready_i_5_22[2] = ready_o_6_22[1];
    data_i_5_22[0] = data_i[5][22];
    valid_i_5_22[0] = valid_i[5][22];
    ready_i_5_22[0] = ready_i[5][22];
end


/*Router 5,23*/    
merge_router #(
    .input_mask                     (input_mask_5_23),
    .output_sel                     (output_sel_5_23)
)router235(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_5_23),
    .valid_i                        (valid_i_5_23),
    .ready_o                        (ready_o_5_23),
    .data_o                         (data_o_5_23),
    .valid_o                        (valid_o_5_23),
    .ready_i                        (ready_i_5_23)
);


always@(*) begin
    data_i_5_23[3] = data_o_5_22[4];
    valid_i_5_23[3] = valid_o_5_22[4];
    ready_i_5_23[3] = ready_o_5_22[4];
    data_i_5_23[4] = data_o_5_24[3];
    valid_i_5_23[4] = valid_o_5_24[3];
    ready_i_5_23[4] = ready_o_5_24[3];
    data_i_5_23[1] = data_o_4_23[2];
    valid_i_5_23[1] = valid_o_4_23[2];
    ready_i_5_23[1] = ready_o_4_23[2];
    data_i_5_23[2] = data_o_6_23[1];
    valid_i_5_23[2] = valid_o_6_23[1];
    ready_i_5_23[2] = ready_o_6_23[1];
    data_i_5_23[0] = data_i[5][23];
    valid_i_5_23[0] = valid_i[5][23];
    ready_i_5_23[0] = ready_i[5][23];
end


/*Router 5,24*/    
merge_router #(
    .input_mask                     (input_mask_5_24),
    .output_sel                     (output_sel_5_24)
)router245(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_5_24),
    .valid_i                        (valid_i_5_24),
    .ready_o                        (ready_o_5_24),
    .data_o                         (data_o_5_24),
    .valid_o                        (valid_o_5_24),
    .ready_i                        (ready_i_5_24)
);


always@(*) begin
    data_i_5_24[3] = data_o_5_23[4];
    valid_i_5_24[3] = valid_o_5_23[4];
    ready_i_5_24[3] = ready_o_5_23[4];
    data_i_5_24[1] = data_o_4_24[2];
    valid_i_5_24[1] = valid_o_4_24[2];
    ready_i_5_24[1] = ready_o_4_24[2];
    data_i_5_24[2] = data_o_6_24[1];
    valid_i_5_24[2] = valid_o_6_24[1];
    ready_i_5_24[2] = ready_o_6_24[1];
    data_i_5_24[0] = data_i[5][24];
    valid_i_5_24[0] = valid_i[5][24];
    ready_i_5_24[0] = ready_i[5][24];
end


/*Router 6,0*/    
merge_router #(
    .input_mask                     (input_mask_6_0),
    .output_sel                     (output_sel_6_0)
)router6(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_6_0),
    .valid_i                        (valid_i_6_0),
    .ready_o                        (ready_o_6_0),
    .data_o                         (data_o_6_0),
    .valid_o                        (valid_o_6_0),
    .ready_i                        (ready_i_6_0)
);


always@(*) begin
    data_i_6_0[4] = data_o_6_1[3];
    valid_i_6_0[4] = valid_o_6_1[3];
    ready_i_6_0[4] = ready_o_6_1[3];
    data_i_6_0[1] = data_o_5_0[2];
    valid_i_6_0[1] = valid_o_5_0[2];
    ready_i_6_0[1] = ready_o_5_0[2];
    data_i_6_0[2] = data_o_7_0[1];
    valid_i_6_0[2] = valid_o_7_0[1];
    ready_i_6_0[2] = ready_o_7_0[1];
    data_i_6_0[0] = data_i[6][0];
    valid_i_6_0[0] = valid_i[6][0];
    ready_i_6_0[0] = ready_i[6][0];
end


/*Router 6,1*/    
merge_router #(
    .input_mask                     (input_mask_6_1),
    .output_sel                     (output_sel_6_1)
)router16(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_6_1),
    .valid_i                        (valid_i_6_1),
    .ready_o                        (ready_o_6_1),
    .data_o                         (data_o_6_1),
    .valid_o                        (valid_o_6_1),
    .ready_i                        (ready_i_6_1)
);


always@(*) begin
    data_i_6_1[3] = data_o_6_0[4];
    valid_i_6_1[3] = valid_o_6_0[4];
    ready_i_6_1[3] = ready_o_6_0[4];
    data_i_6_1[4] = data_o_6_2[3];
    valid_i_6_1[4] = valid_o_6_2[3];
    ready_i_6_1[4] = ready_o_6_2[3];
    data_i_6_1[1] = data_o_5_1[2];
    valid_i_6_1[1] = valid_o_5_1[2];
    ready_i_6_1[1] = ready_o_5_1[2];
    data_i_6_1[2] = data_o_7_1[1];
    valid_i_6_1[2] = valid_o_7_1[1];
    ready_i_6_1[2] = ready_o_7_1[1];
    data_i_6_1[0] = data_i[6][1];
    valid_i_6_1[0] = valid_i[6][1];
    ready_i_6_1[0] = ready_i[6][1];
end


/*Router 6,2*/    
merge_router #(
    .input_mask                     (input_mask_6_2),
    .output_sel                     (output_sel_6_2)
)router26(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_6_2),
    .valid_i                        (valid_i_6_2),
    .ready_o                        (ready_o_6_2),
    .data_o                         (data_o_6_2),
    .valid_o                        (valid_o_6_2),
    .ready_i                        (ready_i_6_2)
);


always@(*) begin
    data_i_6_2[3] = data_o_6_1[4];
    valid_i_6_2[3] = valid_o_6_1[4];
    ready_i_6_2[3] = ready_o_6_1[4];
    data_i_6_2[4] = data_o_6_3[3];
    valid_i_6_2[4] = valid_o_6_3[3];
    ready_i_6_2[4] = ready_o_6_3[3];
    data_i_6_2[1] = data_o_5_2[2];
    valid_i_6_2[1] = valid_o_5_2[2];
    ready_i_6_2[1] = ready_o_5_2[2];
    data_i_6_2[2] = data_o_7_2[1];
    valid_i_6_2[2] = valid_o_7_2[1];
    ready_i_6_2[2] = ready_o_7_2[1];
    data_i_6_2[0] = data_i[6][2];
    valid_i_6_2[0] = valid_i[6][2];
    ready_i_6_2[0] = ready_i[6][2];
end


/*Router 6,3*/    
merge_router #(
    .input_mask                     (input_mask_6_3),
    .output_sel                     (output_sel_6_3)
)router36(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_6_3),
    .valid_i                        (valid_i_6_3),
    .ready_o                        (ready_o_6_3),
    .data_o                         (data_o_6_3),
    .valid_o                        (valid_o_6_3),
    .ready_i                        (ready_i_6_3)
);


always@(*) begin
    data_i_6_3[3] = data_o_6_2[4];
    valid_i_6_3[3] = valid_o_6_2[4];
    ready_i_6_3[3] = ready_o_6_2[4];
    data_i_6_3[4] = data_o_6_4[3];
    valid_i_6_3[4] = valid_o_6_4[3];
    ready_i_6_3[4] = ready_o_6_4[3];
    data_i_6_3[1] = data_o_5_3[2];
    valid_i_6_3[1] = valid_o_5_3[2];
    ready_i_6_3[1] = ready_o_5_3[2];
    data_i_6_3[2] = data_o_7_3[1];
    valid_i_6_3[2] = valid_o_7_3[1];
    ready_i_6_3[2] = ready_o_7_3[1];
    data_i_6_3[0] = data_i[6][3];
    valid_i_6_3[0] = valid_i[6][3];
    ready_i_6_3[0] = ready_i[6][3];
end


/*Router 6,4*/    
merge_router #(
    .input_mask                     (input_mask_6_4),
    .output_sel                     (output_sel_6_4)
)router46(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_6_4),
    .valid_i                        (valid_i_6_4),
    .ready_o                        (ready_o_6_4),
    .data_o                         (data_o_6_4),
    .valid_o                        (valid_o_6_4),
    .ready_i                        (ready_i_6_4)
);


always@(*) begin
    data_i_6_4[3] = data_o_6_3[4];
    valid_i_6_4[3] = valid_o_6_3[4];
    ready_i_6_4[3] = ready_o_6_3[4];
    data_i_6_4[4] = data_o_6_5[3];
    valid_i_6_4[4] = valid_o_6_5[3];
    ready_i_6_4[4] = ready_o_6_5[3];
    data_i_6_4[1] = data_o_5_4[2];
    valid_i_6_4[1] = valid_o_5_4[2];
    ready_i_6_4[1] = ready_o_5_4[2];
    data_i_6_4[2] = data_o_7_4[1];
    valid_i_6_4[2] = valid_o_7_4[1];
    ready_i_6_4[2] = ready_o_7_4[1];
    data_i_6_4[0] = data_i[6][4];
    valid_i_6_4[0] = valid_i[6][4];
    ready_i_6_4[0] = ready_i[6][4];
end


/*Router 6,5*/    
merge_router #(
    .input_mask                     (input_mask_6_5),
    .output_sel                     (output_sel_6_5)
)router56(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_6_5),
    .valid_i                        (valid_i_6_5),
    .ready_o                        (ready_o_6_5),
    .data_o                         (data_o_6_5),
    .valid_o                        (valid_o_6_5),
    .ready_i                        (ready_i_6_5)
);


always@(*) begin
    data_i_6_5[3] = data_o_6_4[4];
    valid_i_6_5[3] = valid_o_6_4[4];
    ready_i_6_5[3] = ready_o_6_4[4];
    data_i_6_5[4] = data_o_6_6[3];
    valid_i_6_5[4] = valid_o_6_6[3];
    ready_i_6_5[4] = ready_o_6_6[3];
    data_i_6_5[1] = data_o_5_5[2];
    valid_i_6_5[1] = valid_o_5_5[2];
    ready_i_6_5[1] = ready_o_5_5[2];
    data_i_6_5[2] = data_o_7_5[1];
    valid_i_6_5[2] = valid_o_7_5[1];
    ready_i_6_5[2] = ready_o_7_5[1];
    data_i_6_5[0] = data_i[6][5];
    valid_i_6_5[0] = valid_i[6][5];
    ready_i_6_5[0] = ready_i[6][5];
end


/*Router 6,6*/    
merge_router #(
    .input_mask                     (input_mask_6_6),
    .output_sel                     (output_sel_6_6)
)router66(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_6_6),
    .valid_i                        (valid_i_6_6),
    .ready_o                        (ready_o_6_6),
    .data_o                         (data_o_6_6),
    .valid_o                        (valid_o_6_6),
    .ready_i                        (ready_i_6_6)
);


always@(*) begin
    data_i_6_6[3] = data_o_6_5[4];
    valid_i_6_6[3] = valid_o_6_5[4];
    ready_i_6_6[3] = ready_o_6_5[4];
    data_i_6_6[4] = data_o_6_7[3];
    valid_i_6_6[4] = valid_o_6_7[3];
    ready_i_6_6[4] = ready_o_6_7[3];
    data_i_6_6[1] = data_o_5_6[2];
    valid_i_6_6[1] = valid_o_5_6[2];
    ready_i_6_6[1] = ready_o_5_6[2];
    data_i_6_6[2] = data_o_7_6[1];
    valid_i_6_6[2] = valid_o_7_6[1];
    ready_i_6_6[2] = ready_o_7_6[1];
    data_i_6_6[0] = data_i[6][6];
    valid_i_6_6[0] = valid_i[6][6];
    ready_i_6_6[0] = ready_i[6][6];
end


/*Router 6,7*/    
merge_router #(
    .input_mask                     (input_mask_6_7),
    .output_sel                     (output_sel_6_7)
)router76(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_6_7),
    .valid_i                        (valid_i_6_7),
    .ready_o                        (ready_o_6_7),
    .data_o                         (data_o_6_7),
    .valid_o                        (valid_o_6_7),
    .ready_i                        (ready_i_6_7)
);


always@(*) begin
    data_i_6_7[3] = data_o_6_6[4];
    valid_i_6_7[3] = valid_o_6_6[4];
    ready_i_6_7[3] = ready_o_6_6[4];
    data_i_6_7[4] = data_o_6_8[3];
    valid_i_6_7[4] = valid_o_6_8[3];
    ready_i_6_7[4] = ready_o_6_8[3];
    data_i_6_7[1] = data_o_5_7[2];
    valid_i_6_7[1] = valid_o_5_7[2];
    ready_i_6_7[1] = ready_o_5_7[2];
    data_i_6_7[2] = data_o_7_7[1];
    valid_i_6_7[2] = valid_o_7_7[1];
    ready_i_6_7[2] = ready_o_7_7[1];
    data_i_6_7[0] = data_i[6][7];
    valid_i_6_7[0] = valid_i[6][7];
    ready_i_6_7[0] = ready_i[6][7];
end


/*Router 6,8*/    
merge_router #(
    .input_mask                     (input_mask_6_8),
    .output_sel                     (output_sel_6_8)
)router86(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_6_8),
    .valid_i                        (valid_i_6_8),
    .ready_o                        (ready_o_6_8),
    .data_o                         (data_o_6_8),
    .valid_o                        (valid_o_6_8),
    .ready_i                        (ready_i_6_8)
);


always@(*) begin
    data_i_6_8[3] = data_o_6_7[4];
    valid_i_6_8[3] = valid_o_6_7[4];
    ready_i_6_8[3] = ready_o_6_7[4];
    data_i_6_8[4] = data_o_6_9[3];
    valid_i_6_8[4] = valid_o_6_9[3];
    ready_i_6_8[4] = ready_o_6_9[3];
    data_i_6_8[1] = data_o_5_8[2];
    valid_i_6_8[1] = valid_o_5_8[2];
    ready_i_6_8[1] = ready_o_5_8[2];
    data_i_6_8[2] = data_o_7_8[1];
    valid_i_6_8[2] = valid_o_7_8[1];
    ready_i_6_8[2] = ready_o_7_8[1];
    data_i_6_8[0] = data_i[6][8];
    valid_i_6_8[0] = valid_i[6][8];
    ready_i_6_8[0] = ready_i[6][8];
end


/*Router 6,9*/    
merge_router #(
    .input_mask                     (input_mask_6_9),
    .output_sel                     (output_sel_6_9)
)router96(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_6_9),
    .valid_i                        (valid_i_6_9),
    .ready_o                        (ready_o_6_9),
    .data_o                         (data_o_6_9),
    .valid_o                        (valid_o_6_9),
    .ready_i                        (ready_i_6_9)
);


always@(*) begin
    data_i_6_9[3] = data_o_6_8[4];
    valid_i_6_9[3] = valid_o_6_8[4];
    ready_i_6_9[3] = ready_o_6_8[4];
    data_i_6_9[4] = data_o_6_10[3];
    valid_i_6_9[4] = valid_o_6_10[3];
    ready_i_6_9[4] = ready_o_6_10[3];
    data_i_6_9[1] = data_o_5_9[2];
    valid_i_6_9[1] = valid_o_5_9[2];
    ready_i_6_9[1] = ready_o_5_9[2];
    data_i_6_9[2] = data_o_7_9[1];
    valid_i_6_9[2] = valid_o_7_9[1];
    ready_i_6_9[2] = ready_o_7_9[1];
    data_i_6_9[0] = data_i[6][9];
    valid_i_6_9[0] = valid_i[6][9];
    ready_i_6_9[0] = ready_i[6][9];
end


/*Router 6,10*/    
merge_router #(
    .input_mask                     (input_mask_6_10),
    .output_sel                     (output_sel_6_10)
)router106(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_6_10),
    .valid_i                        (valid_i_6_10),
    .ready_o                        (ready_o_6_10),
    .data_o                         (data_o_6_10),
    .valid_o                        (valid_o_6_10),
    .ready_i                        (ready_i_6_10)
);


always@(*) begin
    data_i_6_10[3] = data_o_6_9[4];
    valid_i_6_10[3] = valid_o_6_9[4];
    ready_i_6_10[3] = ready_o_6_9[4];
    data_i_6_10[4] = data_o_6_11[3];
    valid_i_6_10[4] = valid_o_6_11[3];
    ready_i_6_10[4] = ready_o_6_11[3];
    data_i_6_10[1] = data_o_5_10[2];
    valid_i_6_10[1] = valid_o_5_10[2];
    ready_i_6_10[1] = ready_o_5_10[2];
    data_i_6_10[2] = data_o_7_10[1];
    valid_i_6_10[2] = valid_o_7_10[1];
    ready_i_6_10[2] = ready_o_7_10[1];
    data_i_6_10[0] = data_i[6][10];
    valid_i_6_10[0] = valid_i[6][10];
    ready_i_6_10[0] = ready_i[6][10];
end


/*Router 6,11*/    
merge_router #(
    .input_mask                     (input_mask_6_11),
    .output_sel                     (output_sel_6_11)
)router116(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_6_11),
    .valid_i                        (valid_i_6_11),
    .ready_o                        (ready_o_6_11),
    .data_o                         (data_o_6_11),
    .valid_o                        (valid_o_6_11),
    .ready_i                        (ready_i_6_11)
);


always@(*) begin
    data_i_6_11[3] = data_o_6_10[4];
    valid_i_6_11[3] = valid_o_6_10[4];
    ready_i_6_11[3] = ready_o_6_10[4];
    data_i_6_11[4] = data_o_6_12[3];
    valid_i_6_11[4] = valid_o_6_12[3];
    ready_i_6_11[4] = ready_o_6_12[3];
    data_i_6_11[1] = data_o_5_11[2];
    valid_i_6_11[1] = valid_o_5_11[2];
    ready_i_6_11[1] = ready_o_5_11[2];
    data_i_6_11[2] = data_o_7_11[1];
    valid_i_6_11[2] = valid_o_7_11[1];
    ready_i_6_11[2] = ready_o_7_11[1];
    data_i_6_11[0] = data_i[6][11];
    valid_i_6_11[0] = valid_i[6][11];
    ready_i_6_11[0] = ready_i[6][11];
end


/*Router 6,12*/    
merge_router #(
    .input_mask                     (input_mask_6_12),
    .output_sel                     (output_sel_6_12)
)router126(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_6_12),
    .valid_i                        (valid_i_6_12),
    .ready_o                        (ready_o_6_12),
    .data_o                         (data_o_6_12),
    .valid_o                        (valid_o_6_12),
    .ready_i                        (ready_i_6_12)
);


always@(*) begin
    data_i_6_12[3] = data_o_6_11[4];
    valid_i_6_12[3] = valid_o_6_11[4];
    ready_i_6_12[3] = ready_o_6_11[4];
    data_i_6_12[4] = data_o_6_13[3];
    valid_i_6_12[4] = valid_o_6_13[3];
    ready_i_6_12[4] = ready_o_6_13[3];
    data_i_6_12[1] = data_o_5_12[2];
    valid_i_6_12[1] = valid_o_5_12[2];
    ready_i_6_12[1] = ready_o_5_12[2];
    data_i_6_12[2] = data_o_7_12[1];
    valid_i_6_12[2] = valid_o_7_12[1];
    ready_i_6_12[2] = ready_o_7_12[1];
    data_i_6_12[0] = data_i[6][12];
    valid_i_6_12[0] = valid_i[6][12];
    ready_i_6_12[0] = ready_i[6][12];
end


/*Router 6,13*/    
merge_router #(
    .input_mask                     (input_mask_6_13),
    .output_sel                     (output_sel_6_13)
)router136(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_6_13),
    .valid_i                        (valid_i_6_13),
    .ready_o                        (ready_o_6_13),
    .data_o                         (data_o_6_13),
    .valid_o                        (valid_o_6_13),
    .ready_i                        (ready_i_6_13)
);


always@(*) begin
    data_i_6_13[3] = data_o_6_12[4];
    valid_i_6_13[3] = valid_o_6_12[4];
    ready_i_6_13[3] = ready_o_6_12[4];
    data_i_6_13[4] = data_o_6_14[3];
    valid_i_6_13[4] = valid_o_6_14[3];
    ready_i_6_13[4] = ready_o_6_14[3];
    data_i_6_13[1] = data_o_5_13[2];
    valid_i_6_13[1] = valid_o_5_13[2];
    ready_i_6_13[1] = ready_o_5_13[2];
    data_i_6_13[2] = data_o_7_13[1];
    valid_i_6_13[2] = valid_o_7_13[1];
    ready_i_6_13[2] = ready_o_7_13[1];
    data_i_6_13[0] = data_i[6][13];
    valid_i_6_13[0] = valid_i[6][13];
    ready_i_6_13[0] = ready_i[6][13];
end


/*Router 6,14*/    
merge_router #(
    .input_mask                     (input_mask_6_14),
    .output_sel                     (output_sel_6_14)
)router146(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_6_14),
    .valid_i                        (valid_i_6_14),
    .ready_o                        (ready_o_6_14),
    .data_o                         (data_o_6_14),
    .valid_o                        (valid_o_6_14),
    .ready_i                        (ready_i_6_14)
);


always@(*) begin
    data_i_6_14[3] = data_o_6_13[4];
    valid_i_6_14[3] = valid_o_6_13[4];
    ready_i_6_14[3] = ready_o_6_13[4];
    data_i_6_14[4] = data_o_6_15[3];
    valid_i_6_14[4] = valid_o_6_15[3];
    ready_i_6_14[4] = ready_o_6_15[3];
    data_i_6_14[1] = data_o_5_14[2];
    valid_i_6_14[1] = valid_o_5_14[2];
    ready_i_6_14[1] = ready_o_5_14[2];
    data_i_6_14[2] = data_o_7_14[1];
    valid_i_6_14[2] = valid_o_7_14[1];
    ready_i_6_14[2] = ready_o_7_14[1];
    data_i_6_14[0] = data_i[6][14];
    valid_i_6_14[0] = valid_i[6][14];
    ready_i_6_14[0] = ready_i[6][14];
end


/*Router 6,15*/    
merge_router #(
    .input_mask                     (input_mask_6_15),
    .output_sel                     (output_sel_6_15)
)router156(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_6_15),
    .valid_i                        (valid_i_6_15),
    .ready_o                        (ready_o_6_15),
    .data_o                         (data_o_6_15),
    .valid_o                        (valid_o_6_15),
    .ready_i                        (ready_i_6_15)
);


always@(*) begin
    data_i_6_15[3] = data_o_6_14[4];
    valid_i_6_15[3] = valid_o_6_14[4];
    ready_i_6_15[3] = ready_o_6_14[4];
    data_i_6_15[4] = data_o_6_16[3];
    valid_i_6_15[4] = valid_o_6_16[3];
    ready_i_6_15[4] = ready_o_6_16[3];
    data_i_6_15[1] = data_o_5_15[2];
    valid_i_6_15[1] = valid_o_5_15[2];
    ready_i_6_15[1] = ready_o_5_15[2];
    data_i_6_15[2] = data_o_7_15[1];
    valid_i_6_15[2] = valid_o_7_15[1];
    ready_i_6_15[2] = ready_o_7_15[1];
    data_i_6_15[0] = data_i[6][15];
    valid_i_6_15[0] = valid_i[6][15];
    ready_i_6_15[0] = ready_i[6][15];
end


/*Router 6,16*/    
merge_router #(
    .input_mask                     (input_mask_6_16),
    .output_sel                     (output_sel_6_16)
)router166(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_6_16),
    .valid_i                        (valid_i_6_16),
    .ready_o                        (ready_o_6_16),
    .data_o                         (data_o_6_16),
    .valid_o                        (valid_o_6_16),
    .ready_i                        (ready_i_6_16)
);


always@(*) begin
    data_i_6_16[3] = data_o_6_15[4];
    valid_i_6_16[3] = valid_o_6_15[4];
    ready_i_6_16[3] = ready_o_6_15[4];
    data_i_6_16[4] = data_o_6_17[3];
    valid_i_6_16[4] = valid_o_6_17[3];
    ready_i_6_16[4] = ready_o_6_17[3];
    data_i_6_16[1] = data_o_5_16[2];
    valid_i_6_16[1] = valid_o_5_16[2];
    ready_i_6_16[1] = ready_o_5_16[2];
    data_i_6_16[2] = data_o_7_16[1];
    valid_i_6_16[2] = valid_o_7_16[1];
    ready_i_6_16[2] = ready_o_7_16[1];
    data_i_6_16[0] = data_i[6][16];
    valid_i_6_16[0] = valid_i[6][16];
    ready_i_6_16[0] = ready_i[6][16];
end


/*Router 6,17*/    
merge_router #(
    .input_mask                     (input_mask_6_17),
    .output_sel                     (output_sel_6_17)
)router176(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_6_17),
    .valid_i                        (valid_i_6_17),
    .ready_o                        (ready_o_6_17),
    .data_o                         (data_o_6_17),
    .valid_o                        (valid_o_6_17),
    .ready_i                        (ready_i_6_17)
);


always@(*) begin
    data_i_6_17[3] = data_o_6_16[4];
    valid_i_6_17[3] = valid_o_6_16[4];
    ready_i_6_17[3] = ready_o_6_16[4];
    data_i_6_17[4] = data_o_6_18[3];
    valid_i_6_17[4] = valid_o_6_18[3];
    ready_i_6_17[4] = ready_o_6_18[3];
    data_i_6_17[1] = data_o_5_17[2];
    valid_i_6_17[1] = valid_o_5_17[2];
    ready_i_6_17[1] = ready_o_5_17[2];
    data_i_6_17[2] = data_o_7_17[1];
    valid_i_6_17[2] = valid_o_7_17[1];
    ready_i_6_17[2] = ready_o_7_17[1];
    data_i_6_17[0] = data_i[6][17];
    valid_i_6_17[0] = valid_i[6][17];
    ready_i_6_17[0] = ready_i[6][17];
end


/*Router 6,18*/    
merge_router #(
    .input_mask                     (input_mask_6_18),
    .output_sel                     (output_sel_6_18)
)router186(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_6_18),
    .valid_i                        (valid_i_6_18),
    .ready_o                        (ready_o_6_18),
    .data_o                         (data_o_6_18),
    .valid_o                        (valid_o_6_18),
    .ready_i                        (ready_i_6_18)
);


always@(*) begin
    data_i_6_18[3] = data_o_6_17[4];
    valid_i_6_18[3] = valid_o_6_17[4];
    ready_i_6_18[3] = ready_o_6_17[4];
    data_i_6_18[4] = data_o_6_19[3];
    valid_i_6_18[4] = valid_o_6_19[3];
    ready_i_6_18[4] = ready_o_6_19[3];
    data_i_6_18[1] = data_o_5_18[2];
    valid_i_6_18[1] = valid_o_5_18[2];
    ready_i_6_18[1] = ready_o_5_18[2];
    data_i_6_18[2] = data_o_7_18[1];
    valid_i_6_18[2] = valid_o_7_18[1];
    ready_i_6_18[2] = ready_o_7_18[1];
    data_i_6_18[0] = data_i[6][18];
    valid_i_6_18[0] = valid_i[6][18];
    ready_i_6_18[0] = ready_i[6][18];
end


/*Router 6,19*/    
merge_router #(
    .input_mask                     (input_mask_6_19),
    .output_sel                     (output_sel_6_19)
)router196(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_6_19),
    .valid_i                        (valid_i_6_19),
    .ready_o                        (ready_o_6_19),
    .data_o                         (data_o_6_19),
    .valid_o                        (valid_o_6_19),
    .ready_i                        (ready_i_6_19)
);


always@(*) begin
    data_i_6_19[3] = data_o_6_18[4];
    valid_i_6_19[3] = valid_o_6_18[4];
    ready_i_6_19[3] = ready_o_6_18[4];
    data_i_6_19[4] = data_o_6_20[3];
    valid_i_6_19[4] = valid_o_6_20[3];
    ready_i_6_19[4] = ready_o_6_20[3];
    data_i_6_19[1] = data_o_5_19[2];
    valid_i_6_19[1] = valid_o_5_19[2];
    ready_i_6_19[1] = ready_o_5_19[2];
    data_i_6_19[2] = data_o_7_19[1];
    valid_i_6_19[2] = valid_o_7_19[1];
    ready_i_6_19[2] = ready_o_7_19[1];
    data_i_6_19[0] = data_i[6][19];
    valid_i_6_19[0] = valid_i[6][19];
    ready_i_6_19[0] = ready_i[6][19];
end


/*Router 6,20*/    
merge_router #(
    .input_mask                     (input_mask_6_20),
    .output_sel                     (output_sel_6_20)
)router206(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_6_20),
    .valid_i                        (valid_i_6_20),
    .ready_o                        (ready_o_6_20),
    .data_o                         (data_o_6_20),
    .valid_o                        (valid_o_6_20),
    .ready_i                        (ready_i_6_20)
);


always@(*) begin
    data_i_6_20[3] = data_o_6_19[4];
    valid_i_6_20[3] = valid_o_6_19[4];
    ready_i_6_20[3] = ready_o_6_19[4];
    data_i_6_20[4] = data_o_6_21[3];
    valid_i_6_20[4] = valid_o_6_21[3];
    ready_i_6_20[4] = ready_o_6_21[3];
    data_i_6_20[1] = data_o_5_20[2];
    valid_i_6_20[1] = valid_o_5_20[2];
    ready_i_6_20[1] = ready_o_5_20[2];
    data_i_6_20[2] = data_o_7_20[1];
    valid_i_6_20[2] = valid_o_7_20[1];
    ready_i_6_20[2] = ready_o_7_20[1];
    data_i_6_20[0] = data_i[6][20];
    valid_i_6_20[0] = valid_i[6][20];
    ready_i_6_20[0] = ready_i[6][20];
end


/*Router 6,21*/    
merge_router #(
    .input_mask                     (input_mask_6_21),
    .output_sel                     (output_sel_6_21)
)router216(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_6_21),
    .valid_i                        (valid_i_6_21),
    .ready_o                        (ready_o_6_21),
    .data_o                         (data_o_6_21),
    .valid_o                        (valid_o_6_21),
    .ready_i                        (ready_i_6_21)
);


always@(*) begin
    data_i_6_21[3] = data_o_6_20[4];
    valid_i_6_21[3] = valid_o_6_20[4];
    ready_i_6_21[3] = ready_o_6_20[4];
    data_i_6_21[4] = data_o_6_22[3];
    valid_i_6_21[4] = valid_o_6_22[3];
    ready_i_6_21[4] = ready_o_6_22[3];
    data_i_6_21[1] = data_o_5_21[2];
    valid_i_6_21[1] = valid_o_5_21[2];
    ready_i_6_21[1] = ready_o_5_21[2];
    data_i_6_21[2] = data_o_7_21[1];
    valid_i_6_21[2] = valid_o_7_21[1];
    ready_i_6_21[2] = ready_o_7_21[1];
    data_i_6_21[0] = data_i[6][21];
    valid_i_6_21[0] = valid_i[6][21];
    ready_i_6_21[0] = ready_i[6][21];
end


/*Router 6,22*/    
merge_router #(
    .input_mask                     (input_mask_6_22),
    .output_sel                     (output_sel_6_22)
)router226(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_6_22),
    .valid_i                        (valid_i_6_22),
    .ready_o                        (ready_o_6_22),
    .data_o                         (data_o_6_22),
    .valid_o                        (valid_o_6_22),
    .ready_i                        (ready_i_6_22)
);


always@(*) begin
    data_i_6_22[3] = data_o_6_21[4];
    valid_i_6_22[3] = valid_o_6_21[4];
    ready_i_6_22[3] = ready_o_6_21[4];
    data_i_6_22[4] = data_o_6_23[3];
    valid_i_6_22[4] = valid_o_6_23[3];
    ready_i_6_22[4] = ready_o_6_23[3];
    data_i_6_22[1] = data_o_5_22[2];
    valid_i_6_22[1] = valid_o_5_22[2];
    ready_i_6_22[1] = ready_o_5_22[2];
    data_i_6_22[2] = data_o_7_22[1];
    valid_i_6_22[2] = valid_o_7_22[1];
    ready_i_6_22[2] = ready_o_7_22[1];
    data_i_6_22[0] = data_i[6][22];
    valid_i_6_22[0] = valid_i[6][22];
    ready_i_6_22[0] = ready_i[6][22];
end


/*Router 6,23*/    
merge_router #(
    .input_mask                     (input_mask_6_23),
    .output_sel                     (output_sel_6_23)
)router236(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_6_23),
    .valid_i                        (valid_i_6_23),
    .ready_o                        (ready_o_6_23),
    .data_o                         (data_o_6_23),
    .valid_o                        (valid_o_6_23),
    .ready_i                        (ready_i_6_23)
);


always@(*) begin
    data_i_6_23[3] = data_o_6_22[4];
    valid_i_6_23[3] = valid_o_6_22[4];
    ready_i_6_23[3] = ready_o_6_22[4];
    data_i_6_23[4] = data_o_6_24[3];
    valid_i_6_23[4] = valid_o_6_24[3];
    ready_i_6_23[4] = ready_o_6_24[3];
    data_i_6_23[1] = data_o_5_23[2];
    valid_i_6_23[1] = valid_o_5_23[2];
    ready_i_6_23[1] = ready_o_5_23[2];
    data_i_6_23[2] = data_o_7_23[1];
    valid_i_6_23[2] = valid_o_7_23[1];
    ready_i_6_23[2] = ready_o_7_23[1];
    data_i_6_23[0] = data_i[6][23];
    valid_i_6_23[0] = valid_i[6][23];
    ready_i_6_23[0] = ready_i[6][23];
end


/*Router 6,24*/    
merge_router #(
    .input_mask                     (input_mask_6_24),
    .output_sel                     (output_sel_6_24)
)router246(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_6_24),
    .valid_i                        (valid_i_6_24),
    .ready_o                        (ready_o_6_24),
    .data_o                         (data_o_6_24),
    .valid_o                        (valid_o_6_24),
    .ready_i                        (ready_i_6_24)
);


always@(*) begin
    data_i_6_24[3] = data_o_6_23[4];
    valid_i_6_24[3] = valid_o_6_23[4];
    ready_i_6_24[3] = ready_o_6_23[4];
    data_i_6_24[1] = data_o_5_24[2];
    valid_i_6_24[1] = valid_o_5_24[2];
    ready_i_6_24[1] = ready_o_5_24[2];
    data_i_6_24[2] = data_o_7_24[1];
    valid_i_6_24[2] = valid_o_7_24[1];
    ready_i_6_24[2] = ready_o_7_24[1];
    data_i_6_24[0] = data_i[6][24];
    valid_i_6_24[0] = valid_i[6][24];
    ready_i_6_24[0] = ready_i[6][24];
end


/*Router 7,0*/    
merge_router #(
    .input_mask                     (input_mask_7_0),
    .output_sel                     (output_sel_7_0)
)router7(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_7_0),
    .valid_i                        (valid_i_7_0),
    .ready_o                        (ready_o_7_0),
    .data_o                         (data_o_7_0),
    .valid_o                        (valid_o_7_0),
    .ready_i                        (ready_i_7_0)
);


always@(*) begin
    data_i_7_0[4] = data_o_7_1[3];
    valid_i_7_0[4] = valid_o_7_1[3];
    ready_i_7_0[4] = ready_o_7_1[3];
    data_i_7_0[1] = data_o_6_0[2];
    valid_i_7_0[1] = valid_o_6_0[2];
    ready_i_7_0[1] = ready_o_6_0[2];
    data_i_7_0[2] = data_o_8_0[1];
    valid_i_7_0[2] = valid_o_8_0[1];
    ready_i_7_0[2] = ready_o_8_0[1];
    data_i_7_0[0] = data_i[7][0];
    valid_i_7_0[0] = valid_i[7][0];
    ready_i_7_0[0] = ready_i[7][0];
end


/*Router 7,1*/    
merge_router #(
    .input_mask                     (input_mask_7_1),
    .output_sel                     (output_sel_7_1)
)router17(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_7_1),
    .valid_i                        (valid_i_7_1),
    .ready_o                        (ready_o_7_1),
    .data_o                         (data_o_7_1),
    .valid_o                        (valid_o_7_1),
    .ready_i                        (ready_i_7_1)
);


always@(*) begin
    data_i_7_1[3] = data_o_7_0[4];
    valid_i_7_1[3] = valid_o_7_0[4];
    ready_i_7_1[3] = ready_o_7_0[4];
    data_i_7_1[4] = data_o_7_2[3];
    valid_i_7_1[4] = valid_o_7_2[3];
    ready_i_7_1[4] = ready_o_7_2[3];
    data_i_7_1[1] = data_o_6_1[2];
    valid_i_7_1[1] = valid_o_6_1[2];
    ready_i_7_1[1] = ready_o_6_1[2];
    data_i_7_1[2] = data_o_8_1[1];
    valid_i_7_1[2] = valid_o_8_1[1];
    ready_i_7_1[2] = ready_o_8_1[1];
    data_i_7_1[0] = data_i[7][1];
    valid_i_7_1[0] = valid_i[7][1];
    ready_i_7_1[0] = ready_i[7][1];
end


/*Router 7,2*/    
merge_router #(
    .input_mask                     (input_mask_7_2),
    .output_sel                     (output_sel_7_2)
)router27(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_7_2),
    .valid_i                        (valid_i_7_2),
    .ready_o                        (ready_o_7_2),
    .data_o                         (data_o_7_2),
    .valid_o                        (valid_o_7_2),
    .ready_i                        (ready_i_7_2)
);


always@(*) begin
    data_i_7_2[3] = data_o_7_1[4];
    valid_i_7_2[3] = valid_o_7_1[4];
    ready_i_7_2[3] = ready_o_7_1[4];
    data_i_7_2[4] = data_o_7_3[3];
    valid_i_7_2[4] = valid_o_7_3[3];
    ready_i_7_2[4] = ready_o_7_3[3];
    data_i_7_2[1] = data_o_6_2[2];
    valid_i_7_2[1] = valid_o_6_2[2];
    ready_i_7_2[1] = ready_o_6_2[2];
    data_i_7_2[2] = data_o_8_2[1];
    valid_i_7_2[2] = valid_o_8_2[1];
    ready_i_7_2[2] = ready_o_8_2[1];
    data_i_7_2[0] = data_i[7][2];
    valid_i_7_2[0] = valid_i[7][2];
    ready_i_7_2[0] = ready_i[7][2];
end


/*Router 7,3*/    
merge_router #(
    .input_mask                     (input_mask_7_3),
    .output_sel                     (output_sel_7_3)
)router37(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_7_3),
    .valid_i                        (valid_i_7_3),
    .ready_o                        (ready_o_7_3),
    .data_o                         (data_o_7_3),
    .valid_o                        (valid_o_7_3),
    .ready_i                        (ready_i_7_3)
);


always@(*) begin
    data_i_7_3[3] = data_o_7_2[4];
    valid_i_7_3[3] = valid_o_7_2[4];
    ready_i_7_3[3] = ready_o_7_2[4];
    data_i_7_3[4] = data_o_7_4[3];
    valid_i_7_3[4] = valid_o_7_4[3];
    ready_i_7_3[4] = ready_o_7_4[3];
    data_i_7_3[1] = data_o_6_3[2];
    valid_i_7_3[1] = valid_o_6_3[2];
    ready_i_7_3[1] = ready_o_6_3[2];
    data_i_7_3[2] = data_o_8_3[1];
    valid_i_7_3[2] = valid_o_8_3[1];
    ready_i_7_3[2] = ready_o_8_3[1];
    data_i_7_3[0] = data_i[7][3];
    valid_i_7_3[0] = valid_i[7][3];
    ready_i_7_3[0] = ready_i[7][3];
end


/*Router 7,4*/    
merge_router #(
    .input_mask                     (input_mask_7_4),
    .output_sel                     (output_sel_7_4)
)router47(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_7_4),
    .valid_i                        (valid_i_7_4),
    .ready_o                        (ready_o_7_4),
    .data_o                         (data_o_7_4),
    .valid_o                        (valid_o_7_4),
    .ready_i                        (ready_i_7_4)
);


always@(*) begin
    data_i_7_4[3] = data_o_7_3[4];
    valid_i_7_4[3] = valid_o_7_3[4];
    ready_i_7_4[3] = ready_o_7_3[4];
    data_i_7_4[4] = data_o_7_5[3];
    valid_i_7_4[4] = valid_o_7_5[3];
    ready_i_7_4[4] = ready_o_7_5[3];
    data_i_7_4[1] = data_o_6_4[2];
    valid_i_7_4[1] = valid_o_6_4[2];
    ready_i_7_4[1] = ready_o_6_4[2];
    data_i_7_4[2] = data_o_8_4[1];
    valid_i_7_4[2] = valid_o_8_4[1];
    ready_i_7_4[2] = ready_o_8_4[1];
    data_i_7_4[0] = data_i[7][4];
    valid_i_7_4[0] = valid_i[7][4];
    ready_i_7_4[0] = ready_i[7][4];
end


/*Router 7,5*/    
merge_router #(
    .input_mask                     (input_mask_7_5),
    .output_sel                     (output_sel_7_5)
)router57(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_7_5),
    .valid_i                        (valid_i_7_5),
    .ready_o                        (ready_o_7_5),
    .data_o                         (data_o_7_5),
    .valid_o                        (valid_o_7_5),
    .ready_i                        (ready_i_7_5)
);


always@(*) begin
    data_i_7_5[3] = data_o_7_4[4];
    valid_i_7_5[3] = valid_o_7_4[4];
    ready_i_7_5[3] = ready_o_7_4[4];
    data_i_7_5[4] = data_o_7_6[3];
    valid_i_7_5[4] = valid_o_7_6[3];
    ready_i_7_5[4] = ready_o_7_6[3];
    data_i_7_5[1] = data_o_6_5[2];
    valid_i_7_5[1] = valid_o_6_5[2];
    ready_i_7_5[1] = ready_o_6_5[2];
    data_i_7_5[2] = data_o_8_5[1];
    valid_i_7_5[2] = valid_o_8_5[1];
    ready_i_7_5[2] = ready_o_8_5[1];
    data_i_7_5[0] = data_i[7][5];
    valid_i_7_5[0] = valid_i[7][5];
    ready_i_7_5[0] = ready_i[7][5];
end


/*Router 7,6*/    
merge_router #(
    .input_mask                     (input_mask_7_6),
    .output_sel                     (output_sel_7_6)
)router67(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_7_6),
    .valid_i                        (valid_i_7_6),
    .ready_o                        (ready_o_7_6),
    .data_o                         (data_o_7_6),
    .valid_o                        (valid_o_7_6),
    .ready_i                        (ready_i_7_6)
);


always@(*) begin
    data_i_7_6[3] = data_o_7_5[4];
    valid_i_7_6[3] = valid_o_7_5[4];
    ready_i_7_6[3] = ready_o_7_5[4];
    data_i_7_6[4] = data_o_7_7[3];
    valid_i_7_6[4] = valid_o_7_7[3];
    ready_i_7_6[4] = ready_o_7_7[3];
    data_i_7_6[1] = data_o_6_6[2];
    valid_i_7_6[1] = valid_o_6_6[2];
    ready_i_7_6[1] = ready_o_6_6[2];
    data_i_7_6[2] = data_o_8_6[1];
    valid_i_7_6[2] = valid_o_8_6[1];
    ready_i_7_6[2] = ready_o_8_6[1];
    data_i_7_6[0] = data_i[7][6];
    valid_i_7_6[0] = valid_i[7][6];
    ready_i_7_6[0] = ready_i[7][6];
end


/*Router 7,7*/    
merge_router #(
    .input_mask                     (input_mask_7_7),
    .output_sel                     (output_sel_7_7)
)router77(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_7_7),
    .valid_i                        (valid_i_7_7),
    .ready_o                        (ready_o_7_7),
    .data_o                         (data_o_7_7),
    .valid_o                        (valid_o_7_7),
    .ready_i                        (ready_i_7_7)
);


always@(*) begin
    data_i_7_7[3] = data_o_7_6[4];
    valid_i_7_7[3] = valid_o_7_6[4];
    ready_i_7_7[3] = ready_o_7_6[4];
    data_i_7_7[4] = data_o_7_8[3];
    valid_i_7_7[4] = valid_o_7_8[3];
    ready_i_7_7[4] = ready_o_7_8[3];
    data_i_7_7[1] = data_o_6_7[2];
    valid_i_7_7[1] = valid_o_6_7[2];
    ready_i_7_7[1] = ready_o_6_7[2];
    data_i_7_7[2] = data_o_8_7[1];
    valid_i_7_7[2] = valid_o_8_7[1];
    ready_i_7_7[2] = ready_o_8_7[1];
    data_i_7_7[0] = data_i[7][7];
    valid_i_7_7[0] = valid_i[7][7];
    ready_i_7_7[0] = ready_i[7][7];
end


/*Router 7,8*/    
merge_router #(
    .input_mask                     (input_mask_7_8),
    .output_sel                     (output_sel_7_8)
)router87(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_7_8),
    .valid_i                        (valid_i_7_8),
    .ready_o                        (ready_o_7_8),
    .data_o                         (data_o_7_8),
    .valid_o                        (valid_o_7_8),
    .ready_i                        (ready_i_7_8)
);


always@(*) begin
    data_i_7_8[3] = data_o_7_7[4];
    valid_i_7_8[3] = valid_o_7_7[4];
    ready_i_7_8[3] = ready_o_7_7[4];
    data_i_7_8[4] = data_o_7_9[3];
    valid_i_7_8[4] = valid_o_7_9[3];
    ready_i_7_8[4] = ready_o_7_9[3];
    data_i_7_8[1] = data_o_6_8[2];
    valid_i_7_8[1] = valid_o_6_8[2];
    ready_i_7_8[1] = ready_o_6_8[2];
    data_i_7_8[2] = data_o_8_8[1];
    valid_i_7_8[2] = valid_o_8_8[1];
    ready_i_7_8[2] = ready_o_8_8[1];
    data_i_7_8[0] = data_i[7][8];
    valid_i_7_8[0] = valid_i[7][8];
    ready_i_7_8[0] = ready_i[7][8];
end


/*Router 7,9*/    
merge_router #(
    .input_mask                     (input_mask_7_9),
    .output_sel                     (output_sel_7_9)
)router97(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_7_9),
    .valid_i                        (valid_i_7_9),
    .ready_o                        (ready_o_7_9),
    .data_o                         (data_o_7_9),
    .valid_o                        (valid_o_7_9),
    .ready_i                        (ready_i_7_9)
);


always@(*) begin
    data_i_7_9[3] = data_o_7_8[4];
    valid_i_7_9[3] = valid_o_7_8[4];
    ready_i_7_9[3] = ready_o_7_8[4];
    data_i_7_9[4] = data_o_7_10[3];
    valid_i_7_9[4] = valid_o_7_10[3];
    ready_i_7_9[4] = ready_o_7_10[3];
    data_i_7_9[1] = data_o_6_9[2];
    valid_i_7_9[1] = valid_o_6_9[2];
    ready_i_7_9[1] = ready_o_6_9[2];
    data_i_7_9[2] = data_o_8_9[1];
    valid_i_7_9[2] = valid_o_8_9[1];
    ready_i_7_9[2] = ready_o_8_9[1];
    data_i_7_9[0] = data_i[7][9];
    valid_i_7_9[0] = valid_i[7][9];
    ready_i_7_9[0] = ready_i[7][9];
end


/*Router 7,10*/    
merge_router #(
    .input_mask                     (input_mask_7_10),
    .output_sel                     (output_sel_7_10)
)router107(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_7_10),
    .valid_i                        (valid_i_7_10),
    .ready_o                        (ready_o_7_10),
    .data_o                         (data_o_7_10),
    .valid_o                        (valid_o_7_10),
    .ready_i                        (ready_i_7_10)
);


always@(*) begin
    data_i_7_10[3] = data_o_7_9[4];
    valid_i_7_10[3] = valid_o_7_9[4];
    ready_i_7_10[3] = ready_o_7_9[4];
    data_i_7_10[4] = data_o_7_11[3];
    valid_i_7_10[4] = valid_o_7_11[3];
    ready_i_7_10[4] = ready_o_7_11[3];
    data_i_7_10[1] = data_o_6_10[2];
    valid_i_7_10[1] = valid_o_6_10[2];
    ready_i_7_10[1] = ready_o_6_10[2];
    data_i_7_10[2] = data_o_8_10[1];
    valid_i_7_10[2] = valid_o_8_10[1];
    ready_i_7_10[2] = ready_o_8_10[1];
    data_i_7_10[0] = data_i[7][10];
    valid_i_7_10[0] = valid_i[7][10];
    ready_i_7_10[0] = ready_i[7][10];
end


/*Router 7,11*/    
merge_router #(
    .input_mask                     (input_mask_7_11),
    .output_sel                     (output_sel_7_11)
)router117(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_7_11),
    .valid_i                        (valid_i_7_11),
    .ready_o                        (ready_o_7_11),
    .data_o                         (data_o_7_11),
    .valid_o                        (valid_o_7_11),
    .ready_i                        (ready_i_7_11)
);


always@(*) begin
    data_i_7_11[3] = data_o_7_10[4];
    valid_i_7_11[3] = valid_o_7_10[4];
    ready_i_7_11[3] = ready_o_7_10[4];
    data_i_7_11[4] = data_o_7_12[3];
    valid_i_7_11[4] = valid_o_7_12[3];
    ready_i_7_11[4] = ready_o_7_12[3];
    data_i_7_11[1] = data_o_6_11[2];
    valid_i_7_11[1] = valid_o_6_11[2];
    ready_i_7_11[1] = ready_o_6_11[2];
    data_i_7_11[2] = data_o_8_11[1];
    valid_i_7_11[2] = valid_o_8_11[1];
    ready_i_7_11[2] = ready_o_8_11[1];
    data_i_7_11[0] = data_i[7][11];
    valid_i_7_11[0] = valid_i[7][11];
    ready_i_7_11[0] = ready_i[7][11];
end


/*Router 7,12*/    
merge_router #(
    .input_mask                     (input_mask_7_12),
    .output_sel                     (output_sel_7_12)
)router127(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_7_12),
    .valid_i                        (valid_i_7_12),
    .ready_o                        (ready_o_7_12),
    .data_o                         (data_o_7_12),
    .valid_o                        (valid_o_7_12),
    .ready_i                        (ready_i_7_12)
);


always@(*) begin
    data_i_7_12[3] = data_o_7_11[4];
    valid_i_7_12[3] = valid_o_7_11[4];
    ready_i_7_12[3] = ready_o_7_11[4];
    data_i_7_12[4] = data_o_7_13[3];
    valid_i_7_12[4] = valid_o_7_13[3];
    ready_i_7_12[4] = ready_o_7_13[3];
    data_i_7_12[1] = data_o_6_12[2];
    valid_i_7_12[1] = valid_o_6_12[2];
    ready_i_7_12[1] = ready_o_6_12[2];
    data_i_7_12[2] = data_o_8_12[1];
    valid_i_7_12[2] = valid_o_8_12[1];
    ready_i_7_12[2] = ready_o_8_12[1];
    data_i_7_12[0] = data_i[7][12];
    valid_i_7_12[0] = valid_i[7][12];
    ready_i_7_12[0] = ready_i[7][12];
end


/*Router 7,13*/    
merge_router #(
    .input_mask                     (input_mask_7_13),
    .output_sel                     (output_sel_7_13)
)router137(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_7_13),
    .valid_i                        (valid_i_7_13),
    .ready_o                        (ready_o_7_13),
    .data_o                         (data_o_7_13),
    .valid_o                        (valid_o_7_13),
    .ready_i                        (ready_i_7_13)
);


always@(*) begin
    data_i_7_13[3] = data_o_7_12[4];
    valid_i_7_13[3] = valid_o_7_12[4];
    ready_i_7_13[3] = ready_o_7_12[4];
    data_i_7_13[4] = data_o_7_14[3];
    valid_i_7_13[4] = valid_o_7_14[3];
    ready_i_7_13[4] = ready_o_7_14[3];
    data_i_7_13[1] = data_o_6_13[2];
    valid_i_7_13[1] = valid_o_6_13[2];
    ready_i_7_13[1] = ready_o_6_13[2];
    data_i_7_13[2] = data_o_8_13[1];
    valid_i_7_13[2] = valid_o_8_13[1];
    ready_i_7_13[2] = ready_o_8_13[1];
    data_i_7_13[0] = data_i[7][13];
    valid_i_7_13[0] = valid_i[7][13];
    ready_i_7_13[0] = ready_i[7][13];
end


/*Router 7,14*/    
merge_router #(
    .input_mask                     (input_mask_7_14),
    .output_sel                     (output_sel_7_14)
)router147(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_7_14),
    .valid_i                        (valid_i_7_14),
    .ready_o                        (ready_o_7_14),
    .data_o                         (data_o_7_14),
    .valid_o                        (valid_o_7_14),
    .ready_i                        (ready_i_7_14)
);


always@(*) begin
    data_i_7_14[3] = data_o_7_13[4];
    valid_i_7_14[3] = valid_o_7_13[4];
    ready_i_7_14[3] = ready_o_7_13[4];
    data_i_7_14[4] = data_o_7_15[3];
    valid_i_7_14[4] = valid_o_7_15[3];
    ready_i_7_14[4] = ready_o_7_15[3];
    data_i_7_14[1] = data_o_6_14[2];
    valid_i_7_14[1] = valid_o_6_14[2];
    ready_i_7_14[1] = ready_o_6_14[2];
    data_i_7_14[2] = data_o_8_14[1];
    valid_i_7_14[2] = valid_o_8_14[1];
    ready_i_7_14[2] = ready_o_8_14[1];
    data_i_7_14[0] = data_i[7][14];
    valid_i_7_14[0] = valid_i[7][14];
    ready_i_7_14[0] = ready_i[7][14];
end


/*Router 7,15*/    
merge_router #(
    .input_mask                     (input_mask_7_15),
    .output_sel                     (output_sel_7_15)
)router157(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_7_15),
    .valid_i                        (valid_i_7_15),
    .ready_o                        (ready_o_7_15),
    .data_o                         (data_o_7_15),
    .valid_o                        (valid_o_7_15),
    .ready_i                        (ready_i_7_15)
);


always@(*) begin
    data_i_7_15[3] = data_o_7_14[4];
    valid_i_7_15[3] = valid_o_7_14[4];
    ready_i_7_15[3] = ready_o_7_14[4];
    data_i_7_15[4] = data_o_7_16[3];
    valid_i_7_15[4] = valid_o_7_16[3];
    ready_i_7_15[4] = ready_o_7_16[3];
    data_i_7_15[1] = data_o_6_15[2];
    valid_i_7_15[1] = valid_o_6_15[2];
    ready_i_7_15[1] = ready_o_6_15[2];
    data_i_7_15[2] = data_o_8_15[1];
    valid_i_7_15[2] = valid_o_8_15[1];
    ready_i_7_15[2] = ready_o_8_15[1];
    data_i_7_15[0] = data_i[7][15];
    valid_i_7_15[0] = valid_i[7][15];
    ready_i_7_15[0] = ready_i[7][15];
end


/*Router 7,16*/    
merge_router #(
    .input_mask                     (input_mask_7_16),
    .output_sel                     (output_sel_7_16)
)router167(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_7_16),
    .valid_i                        (valid_i_7_16),
    .ready_o                        (ready_o_7_16),
    .data_o                         (data_o_7_16),
    .valid_o                        (valid_o_7_16),
    .ready_i                        (ready_i_7_16)
);


always@(*) begin
    data_i_7_16[3] = data_o_7_15[4];
    valid_i_7_16[3] = valid_o_7_15[4];
    ready_i_7_16[3] = ready_o_7_15[4];
    data_i_7_16[4] = data_o_7_17[3];
    valid_i_7_16[4] = valid_o_7_17[3];
    ready_i_7_16[4] = ready_o_7_17[3];
    data_i_7_16[1] = data_o_6_16[2];
    valid_i_7_16[1] = valid_o_6_16[2];
    ready_i_7_16[1] = ready_o_6_16[2];
    data_i_7_16[2] = data_o_8_16[1];
    valid_i_7_16[2] = valid_o_8_16[1];
    ready_i_7_16[2] = ready_o_8_16[1];
    data_i_7_16[0] = data_i[7][16];
    valid_i_7_16[0] = valid_i[7][16];
    ready_i_7_16[0] = ready_i[7][16];
end


/*Router 7,17*/    
merge_router #(
    .input_mask                     (input_mask_7_17),
    .output_sel                     (output_sel_7_17)
)router177(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_7_17),
    .valid_i                        (valid_i_7_17),
    .ready_o                        (ready_o_7_17),
    .data_o                         (data_o_7_17),
    .valid_o                        (valid_o_7_17),
    .ready_i                        (ready_i_7_17)
);


always@(*) begin
    data_i_7_17[3] = data_o_7_16[4];
    valid_i_7_17[3] = valid_o_7_16[4];
    ready_i_7_17[3] = ready_o_7_16[4];
    data_i_7_17[4] = data_o_7_18[3];
    valid_i_7_17[4] = valid_o_7_18[3];
    ready_i_7_17[4] = ready_o_7_18[3];
    data_i_7_17[1] = data_o_6_17[2];
    valid_i_7_17[1] = valid_o_6_17[2];
    ready_i_7_17[1] = ready_o_6_17[2];
    data_i_7_17[2] = data_o_8_17[1];
    valid_i_7_17[2] = valid_o_8_17[1];
    ready_i_7_17[2] = ready_o_8_17[1];
    data_i_7_17[0] = data_i[7][17];
    valid_i_7_17[0] = valid_i[7][17];
    ready_i_7_17[0] = ready_i[7][17];
end


/*Router 7,18*/    
merge_router #(
    .input_mask                     (input_mask_7_18),
    .output_sel                     (output_sel_7_18)
)router187(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_7_18),
    .valid_i                        (valid_i_7_18),
    .ready_o                        (ready_o_7_18),
    .data_o                         (data_o_7_18),
    .valid_o                        (valid_o_7_18),
    .ready_i                        (ready_i_7_18)
);


always@(*) begin
    data_i_7_18[3] = data_o_7_17[4];
    valid_i_7_18[3] = valid_o_7_17[4];
    ready_i_7_18[3] = ready_o_7_17[4];
    data_i_7_18[4] = data_o_7_19[3];
    valid_i_7_18[4] = valid_o_7_19[3];
    ready_i_7_18[4] = ready_o_7_19[3];
    data_i_7_18[1] = data_o_6_18[2];
    valid_i_7_18[1] = valid_o_6_18[2];
    ready_i_7_18[1] = ready_o_6_18[2];
    data_i_7_18[2] = data_o_8_18[1];
    valid_i_7_18[2] = valid_o_8_18[1];
    ready_i_7_18[2] = ready_o_8_18[1];
    data_i_7_18[0] = data_i[7][18];
    valid_i_7_18[0] = valid_i[7][18];
    ready_i_7_18[0] = ready_i[7][18];
end


/*Router 7,19*/    
merge_router #(
    .input_mask                     (input_mask_7_19),
    .output_sel                     (output_sel_7_19)
)router197(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_7_19),
    .valid_i                        (valid_i_7_19),
    .ready_o                        (ready_o_7_19),
    .data_o                         (data_o_7_19),
    .valid_o                        (valid_o_7_19),
    .ready_i                        (ready_i_7_19)
);


always@(*) begin
    data_i_7_19[3] = data_o_7_18[4];
    valid_i_7_19[3] = valid_o_7_18[4];
    ready_i_7_19[3] = ready_o_7_18[4];
    data_i_7_19[4] = data_o_7_20[3];
    valid_i_7_19[4] = valid_o_7_20[3];
    ready_i_7_19[4] = ready_o_7_20[3];
    data_i_7_19[1] = data_o_6_19[2];
    valid_i_7_19[1] = valid_o_6_19[2];
    ready_i_7_19[1] = ready_o_6_19[2];
    data_i_7_19[2] = data_o_8_19[1];
    valid_i_7_19[2] = valid_o_8_19[1];
    ready_i_7_19[2] = ready_o_8_19[1];
    data_i_7_19[0] = data_i[7][19];
    valid_i_7_19[0] = valid_i[7][19];
    ready_i_7_19[0] = ready_i[7][19];
end


/*Router 7,20*/    
merge_router #(
    .input_mask                     (input_mask_7_20),
    .output_sel                     (output_sel_7_20)
)router207(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_7_20),
    .valid_i                        (valid_i_7_20),
    .ready_o                        (ready_o_7_20),
    .data_o                         (data_o_7_20),
    .valid_o                        (valid_o_7_20),
    .ready_i                        (ready_i_7_20)
);


always@(*) begin
    data_i_7_20[3] = data_o_7_19[4];
    valid_i_7_20[3] = valid_o_7_19[4];
    ready_i_7_20[3] = ready_o_7_19[4];
    data_i_7_20[4] = data_o_7_21[3];
    valid_i_7_20[4] = valid_o_7_21[3];
    ready_i_7_20[4] = ready_o_7_21[3];
    data_i_7_20[1] = data_o_6_20[2];
    valid_i_7_20[1] = valid_o_6_20[2];
    ready_i_7_20[1] = ready_o_6_20[2];
    data_i_7_20[2] = data_o_8_20[1];
    valid_i_7_20[2] = valid_o_8_20[1];
    ready_i_7_20[2] = ready_o_8_20[1];
    data_i_7_20[0] = data_i[7][20];
    valid_i_7_20[0] = valid_i[7][20];
    ready_i_7_20[0] = ready_i[7][20];
end


/*Router 7,21*/    
merge_router #(
    .input_mask                     (input_mask_7_21),
    .output_sel                     (output_sel_7_21)
)router217(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_7_21),
    .valid_i                        (valid_i_7_21),
    .ready_o                        (ready_o_7_21),
    .data_o                         (data_o_7_21),
    .valid_o                        (valid_o_7_21),
    .ready_i                        (ready_i_7_21)
);


always@(*) begin
    data_i_7_21[3] = data_o_7_20[4];
    valid_i_7_21[3] = valid_o_7_20[4];
    ready_i_7_21[3] = ready_o_7_20[4];
    data_i_7_21[4] = data_o_7_22[3];
    valid_i_7_21[4] = valid_o_7_22[3];
    ready_i_7_21[4] = ready_o_7_22[3];
    data_i_7_21[1] = data_o_6_21[2];
    valid_i_7_21[1] = valid_o_6_21[2];
    ready_i_7_21[1] = ready_o_6_21[2];
    data_i_7_21[2] = data_o_8_21[1];
    valid_i_7_21[2] = valid_o_8_21[1];
    ready_i_7_21[2] = ready_o_8_21[1];
    data_i_7_21[0] = data_i[7][21];
    valid_i_7_21[0] = valid_i[7][21];
    ready_i_7_21[0] = ready_i[7][21];
end


/*Router 7,22*/    
merge_router #(
    .input_mask                     (input_mask_7_22),
    .output_sel                     (output_sel_7_22)
)router227(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_7_22),
    .valid_i                        (valid_i_7_22),
    .ready_o                        (ready_o_7_22),
    .data_o                         (data_o_7_22),
    .valid_o                        (valid_o_7_22),
    .ready_i                        (ready_i_7_22)
);


always@(*) begin
    data_i_7_22[3] = data_o_7_21[4];
    valid_i_7_22[3] = valid_o_7_21[4];
    ready_i_7_22[3] = ready_o_7_21[4];
    data_i_7_22[4] = data_o_7_23[3];
    valid_i_7_22[4] = valid_o_7_23[3];
    ready_i_7_22[4] = ready_o_7_23[3];
    data_i_7_22[1] = data_o_6_22[2];
    valid_i_7_22[1] = valid_o_6_22[2];
    ready_i_7_22[1] = ready_o_6_22[2];
    data_i_7_22[2] = data_o_8_22[1];
    valid_i_7_22[2] = valid_o_8_22[1];
    ready_i_7_22[2] = ready_o_8_22[1];
    data_i_7_22[0] = data_i[7][22];
    valid_i_7_22[0] = valid_i[7][22];
    ready_i_7_22[0] = ready_i[7][22];
end


/*Router 7,23*/    
merge_router #(
    .input_mask                     (input_mask_7_23),
    .output_sel                     (output_sel_7_23)
)router237(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_7_23),
    .valid_i                        (valid_i_7_23),
    .ready_o                        (ready_o_7_23),
    .data_o                         (data_o_7_23),
    .valid_o                        (valid_o_7_23),
    .ready_i                        (ready_i_7_23)
);


always@(*) begin
    data_i_7_23[3] = data_o_7_22[4];
    valid_i_7_23[3] = valid_o_7_22[4];
    ready_i_7_23[3] = ready_o_7_22[4];
    data_i_7_23[4] = data_o_7_24[3];
    valid_i_7_23[4] = valid_o_7_24[3];
    ready_i_7_23[4] = ready_o_7_24[3];
    data_i_7_23[1] = data_o_6_23[2];
    valid_i_7_23[1] = valid_o_6_23[2];
    ready_i_7_23[1] = ready_o_6_23[2];
    data_i_7_23[2] = data_o_8_23[1];
    valid_i_7_23[2] = valid_o_8_23[1];
    ready_i_7_23[2] = ready_o_8_23[1];
    data_i_7_23[0] = data_i[7][23];
    valid_i_7_23[0] = valid_i[7][23];
    ready_i_7_23[0] = ready_i[7][23];
end


/*Router 7,24*/    
merge_router #(
    .input_mask                     (input_mask_7_24),
    .output_sel                     (output_sel_7_24)
)router247(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_7_24),
    .valid_i                        (valid_i_7_24),
    .ready_o                        (ready_o_7_24),
    .data_o                         (data_o_7_24),
    .valid_o                        (valid_o_7_24),
    .ready_i                        (ready_i_7_24)
);


always@(*) begin
    data_i_7_24[3] = data_o_7_23[4];
    valid_i_7_24[3] = valid_o_7_23[4];
    ready_i_7_24[3] = ready_o_7_23[4];
    data_i_7_24[1] = data_o_6_24[2];
    valid_i_7_24[1] = valid_o_6_24[2];
    ready_i_7_24[1] = ready_o_6_24[2];
    data_i_7_24[2] = data_o_8_24[1];
    valid_i_7_24[2] = valid_o_8_24[1];
    ready_i_7_24[2] = ready_o_8_24[1];
    data_i_7_24[0] = data_i[7][24];
    valid_i_7_24[0] = valid_i[7][24];
    ready_i_7_24[0] = ready_i[7][24];
end


/*Router 8,0*/    
merge_router #(
    .input_mask                     (input_mask_8_0),
    .output_sel                     (output_sel_8_0)
)router8(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_8_0),
    .valid_i                        (valid_i_8_0),
    .ready_o                        (ready_o_8_0),
    .data_o                         (data_o_8_0),
    .valid_o                        (valid_o_8_0),
    .ready_i                        (ready_i_8_0)
);


always@(*) begin
    data_i_8_0[4] = data_o_8_1[3];
    valid_i_8_0[4] = valid_o_8_1[3];
    ready_i_8_0[4] = ready_o_8_1[3];
    data_i_8_0[1] = data_o_7_0[2];
    valid_i_8_0[1] = valid_o_7_0[2];
    ready_i_8_0[1] = ready_o_7_0[2];
    data_i_8_0[2] = data_o_9_0[1];
    valid_i_8_0[2] = valid_o_9_0[1];
    ready_i_8_0[2] = ready_o_9_0[1];
    data_i_8_0[0] = data_i[8][0];
    valid_i_8_0[0] = valid_i[8][0];
    ready_i_8_0[0] = ready_i[8][0];
end


/*Router 8,1*/    
merge_router #(
    .input_mask                     (input_mask_8_1),
    .output_sel                     (output_sel_8_1)
)router18(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_8_1),
    .valid_i                        (valid_i_8_1),
    .ready_o                        (ready_o_8_1),
    .data_o                         (data_o_8_1),
    .valid_o                        (valid_o_8_1),
    .ready_i                        (ready_i_8_1)
);


always@(*) begin
    data_i_8_1[3] = data_o_8_0[4];
    valid_i_8_1[3] = valid_o_8_0[4];
    ready_i_8_1[3] = ready_o_8_0[4];
    data_i_8_1[4] = data_o_8_2[3];
    valid_i_8_1[4] = valid_o_8_2[3];
    ready_i_8_1[4] = ready_o_8_2[3];
    data_i_8_1[1] = data_o_7_1[2];
    valid_i_8_1[1] = valid_o_7_1[2];
    ready_i_8_1[1] = ready_o_7_1[2];
    data_i_8_1[2] = data_o_9_1[1];
    valid_i_8_1[2] = valid_o_9_1[1];
    ready_i_8_1[2] = ready_o_9_1[1];
    data_i_8_1[0] = data_i[8][1];
    valid_i_8_1[0] = valid_i[8][1];
    ready_i_8_1[0] = ready_i[8][1];
end


/*Router 8,2*/    
merge_router #(
    .input_mask                     (input_mask_8_2),
    .output_sel                     (output_sel_8_2)
)router28(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_8_2),
    .valid_i                        (valid_i_8_2),
    .ready_o                        (ready_o_8_2),
    .data_o                         (data_o_8_2),
    .valid_o                        (valid_o_8_2),
    .ready_i                        (ready_i_8_2)
);


always@(*) begin
    data_i_8_2[3] = data_o_8_1[4];
    valid_i_8_2[3] = valid_o_8_1[4];
    ready_i_8_2[3] = ready_o_8_1[4];
    data_i_8_2[4] = data_o_8_3[3];
    valid_i_8_2[4] = valid_o_8_3[3];
    ready_i_8_2[4] = ready_o_8_3[3];
    data_i_8_2[1] = data_o_7_2[2];
    valid_i_8_2[1] = valid_o_7_2[2];
    ready_i_8_2[1] = ready_o_7_2[2];
    data_i_8_2[2] = data_o_9_2[1];
    valid_i_8_2[2] = valid_o_9_2[1];
    ready_i_8_2[2] = ready_o_9_2[1];
    data_i_8_2[0] = data_i[8][2];
    valid_i_8_2[0] = valid_i[8][2];
    ready_i_8_2[0] = ready_i[8][2];
end


/*Router 8,3*/    
merge_router #(
    .input_mask                     (input_mask_8_3),
    .output_sel                     (output_sel_8_3)
)router38(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_8_3),
    .valid_i                        (valid_i_8_3),
    .ready_o                        (ready_o_8_3),
    .data_o                         (data_o_8_3),
    .valid_o                        (valid_o_8_3),
    .ready_i                        (ready_i_8_3)
);


always@(*) begin
    data_i_8_3[3] = data_o_8_2[4];
    valid_i_8_3[3] = valid_o_8_2[4];
    ready_i_8_3[3] = ready_o_8_2[4];
    data_i_8_3[4] = data_o_8_4[3];
    valid_i_8_3[4] = valid_o_8_4[3];
    ready_i_8_3[4] = ready_o_8_4[3];
    data_i_8_3[1] = data_o_7_3[2];
    valid_i_8_3[1] = valid_o_7_3[2];
    ready_i_8_3[1] = ready_o_7_3[2];
    data_i_8_3[2] = data_o_9_3[1];
    valid_i_8_3[2] = valid_o_9_3[1];
    ready_i_8_3[2] = ready_o_9_3[1];
    data_i_8_3[0] = data_i[8][3];
    valid_i_8_3[0] = valid_i[8][3];
    ready_i_8_3[0] = ready_i[8][3];
end


/*Router 8,4*/    
merge_router #(
    .input_mask                     (input_mask_8_4),
    .output_sel                     (output_sel_8_4)
)router48(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_8_4),
    .valid_i                        (valid_i_8_4),
    .ready_o                        (ready_o_8_4),
    .data_o                         (data_o_8_4),
    .valid_o                        (valid_o_8_4),
    .ready_i                        (ready_i_8_4)
);


always@(*) begin
    data_i_8_4[3] = data_o_8_3[4];
    valid_i_8_4[3] = valid_o_8_3[4];
    ready_i_8_4[3] = ready_o_8_3[4];
    data_i_8_4[4] = data_o_8_5[3];
    valid_i_8_4[4] = valid_o_8_5[3];
    ready_i_8_4[4] = ready_o_8_5[3];
    data_i_8_4[1] = data_o_7_4[2];
    valid_i_8_4[1] = valid_o_7_4[2];
    ready_i_8_4[1] = ready_o_7_4[2];
    data_i_8_4[2] = data_o_9_4[1];
    valid_i_8_4[2] = valid_o_9_4[1];
    ready_i_8_4[2] = ready_o_9_4[1];
    data_i_8_4[0] = data_i[8][4];
    valid_i_8_4[0] = valid_i[8][4];
    ready_i_8_4[0] = ready_i[8][4];
end


/*Router 8,5*/    
merge_router #(
    .input_mask                     (input_mask_8_5),
    .output_sel                     (output_sel_8_5)
)router58(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_8_5),
    .valid_i                        (valid_i_8_5),
    .ready_o                        (ready_o_8_5),
    .data_o                         (data_o_8_5),
    .valid_o                        (valid_o_8_5),
    .ready_i                        (ready_i_8_5)
);


always@(*) begin
    data_i_8_5[3] = data_o_8_4[4];
    valid_i_8_5[3] = valid_o_8_4[4];
    ready_i_8_5[3] = ready_o_8_4[4];
    data_i_8_5[4] = data_o_8_6[3];
    valid_i_8_5[4] = valid_o_8_6[3];
    ready_i_8_5[4] = ready_o_8_6[3];
    data_i_8_5[1] = data_o_7_5[2];
    valid_i_8_5[1] = valid_o_7_5[2];
    ready_i_8_5[1] = ready_o_7_5[2];
    data_i_8_5[2] = data_o_9_5[1];
    valid_i_8_5[2] = valid_o_9_5[1];
    ready_i_8_5[2] = ready_o_9_5[1];
    data_i_8_5[0] = data_i[8][5];
    valid_i_8_5[0] = valid_i[8][5];
    ready_i_8_5[0] = ready_i[8][5];
end


/*Router 8,6*/    
merge_router #(
    .input_mask                     (input_mask_8_6),
    .output_sel                     (output_sel_8_6)
)router68(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_8_6),
    .valid_i                        (valid_i_8_6),
    .ready_o                        (ready_o_8_6),
    .data_o                         (data_o_8_6),
    .valid_o                        (valid_o_8_6),
    .ready_i                        (ready_i_8_6)
);


always@(*) begin
    data_i_8_6[3] = data_o_8_5[4];
    valid_i_8_6[3] = valid_o_8_5[4];
    ready_i_8_6[3] = ready_o_8_5[4];
    data_i_8_6[4] = data_o_8_7[3];
    valid_i_8_6[4] = valid_o_8_7[3];
    ready_i_8_6[4] = ready_o_8_7[3];
    data_i_8_6[1] = data_o_7_6[2];
    valid_i_8_6[1] = valid_o_7_6[2];
    ready_i_8_6[1] = ready_o_7_6[2];
    data_i_8_6[2] = data_o_9_6[1];
    valid_i_8_6[2] = valid_o_9_6[1];
    ready_i_8_6[2] = ready_o_9_6[1];
    data_i_8_6[0] = data_i[8][6];
    valid_i_8_6[0] = valid_i[8][6];
    ready_i_8_6[0] = ready_i[8][6];
end


/*Router 8,7*/    
merge_router #(
    .input_mask                     (input_mask_8_7),
    .output_sel                     (output_sel_8_7)
)router78(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_8_7),
    .valid_i                        (valid_i_8_7),
    .ready_o                        (ready_o_8_7),
    .data_o                         (data_o_8_7),
    .valid_o                        (valid_o_8_7),
    .ready_i                        (ready_i_8_7)
);


always@(*) begin
    data_i_8_7[3] = data_o_8_6[4];
    valid_i_8_7[3] = valid_o_8_6[4];
    ready_i_8_7[3] = ready_o_8_6[4];
    data_i_8_7[4] = data_o_8_8[3];
    valid_i_8_7[4] = valid_o_8_8[3];
    ready_i_8_7[4] = ready_o_8_8[3];
    data_i_8_7[1] = data_o_7_7[2];
    valid_i_8_7[1] = valid_o_7_7[2];
    ready_i_8_7[1] = ready_o_7_7[2];
    data_i_8_7[2] = data_o_9_7[1];
    valid_i_8_7[2] = valid_o_9_7[1];
    ready_i_8_7[2] = ready_o_9_7[1];
    data_i_8_7[0] = data_i[8][7];
    valid_i_8_7[0] = valid_i[8][7];
    ready_i_8_7[0] = ready_i[8][7];
end


/*Router 8,8*/    
merge_router #(
    .input_mask                     (input_mask_8_8),
    .output_sel                     (output_sel_8_8)
)router88(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_8_8),
    .valid_i                        (valid_i_8_8),
    .ready_o                        (ready_o_8_8),
    .data_o                         (data_o_8_8),
    .valid_o                        (valid_o_8_8),
    .ready_i                        (ready_i_8_8)
);


always@(*) begin
    data_i_8_8[3] = data_o_8_7[4];
    valid_i_8_8[3] = valid_o_8_7[4];
    ready_i_8_8[3] = ready_o_8_7[4];
    data_i_8_8[4] = data_o_8_9[3];
    valid_i_8_8[4] = valid_o_8_9[3];
    ready_i_8_8[4] = ready_o_8_9[3];
    data_i_8_8[1] = data_o_7_8[2];
    valid_i_8_8[1] = valid_o_7_8[2];
    ready_i_8_8[1] = ready_o_7_8[2];
    data_i_8_8[2] = data_o_9_8[1];
    valid_i_8_8[2] = valid_o_9_8[1];
    ready_i_8_8[2] = ready_o_9_8[1];
    data_i_8_8[0] = data_i[8][8];
    valid_i_8_8[0] = valid_i[8][8];
    ready_i_8_8[0] = ready_i[8][8];
end


/*Router 8,9*/    
merge_router #(
    .input_mask                     (input_mask_8_9),
    .output_sel                     (output_sel_8_9)
)router98(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_8_9),
    .valid_i                        (valid_i_8_9),
    .ready_o                        (ready_o_8_9),
    .data_o                         (data_o_8_9),
    .valid_o                        (valid_o_8_9),
    .ready_i                        (ready_i_8_9)
);


always@(*) begin
    data_i_8_9[3] = data_o_8_8[4];
    valid_i_8_9[3] = valid_o_8_8[4];
    ready_i_8_9[3] = ready_o_8_8[4];
    data_i_8_9[4] = data_o_8_10[3];
    valid_i_8_9[4] = valid_o_8_10[3];
    ready_i_8_9[4] = ready_o_8_10[3];
    data_i_8_9[1] = data_o_7_9[2];
    valid_i_8_9[1] = valid_o_7_9[2];
    ready_i_8_9[1] = ready_o_7_9[2];
    data_i_8_9[2] = data_o_9_9[1];
    valid_i_8_9[2] = valid_o_9_9[1];
    ready_i_8_9[2] = ready_o_9_9[1];
    data_i_8_9[0] = data_i[8][9];
    valid_i_8_9[0] = valid_i[8][9];
    ready_i_8_9[0] = ready_i[8][9];
end


/*Router 8,10*/    
merge_router #(
    .input_mask                     (input_mask_8_10),
    .output_sel                     (output_sel_8_10)
)router108(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_8_10),
    .valid_i                        (valid_i_8_10),
    .ready_o                        (ready_o_8_10),
    .data_o                         (data_o_8_10),
    .valid_o                        (valid_o_8_10),
    .ready_i                        (ready_i_8_10)
);


always@(*) begin
    data_i_8_10[3] = data_o_8_9[4];
    valid_i_8_10[3] = valid_o_8_9[4];
    ready_i_8_10[3] = ready_o_8_9[4];
    data_i_8_10[4] = data_o_8_11[3];
    valid_i_8_10[4] = valid_o_8_11[3];
    ready_i_8_10[4] = ready_o_8_11[3];
    data_i_8_10[1] = data_o_7_10[2];
    valid_i_8_10[1] = valid_o_7_10[2];
    ready_i_8_10[1] = ready_o_7_10[2];
    data_i_8_10[2] = data_o_9_10[1];
    valid_i_8_10[2] = valid_o_9_10[1];
    ready_i_8_10[2] = ready_o_9_10[1];
    data_i_8_10[0] = data_i[8][10];
    valid_i_8_10[0] = valid_i[8][10];
    ready_i_8_10[0] = ready_i[8][10];
end


/*Router 8,11*/    
merge_router #(
    .input_mask                     (input_mask_8_11),
    .output_sel                     (output_sel_8_11)
)router118(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_8_11),
    .valid_i                        (valid_i_8_11),
    .ready_o                        (ready_o_8_11),
    .data_o                         (data_o_8_11),
    .valid_o                        (valid_o_8_11),
    .ready_i                        (ready_i_8_11)
);


always@(*) begin
    data_i_8_11[3] = data_o_8_10[4];
    valid_i_8_11[3] = valid_o_8_10[4];
    ready_i_8_11[3] = ready_o_8_10[4];
    data_i_8_11[4] = data_o_8_12[3];
    valid_i_8_11[4] = valid_o_8_12[3];
    ready_i_8_11[4] = ready_o_8_12[3];
    data_i_8_11[1] = data_o_7_11[2];
    valid_i_8_11[1] = valid_o_7_11[2];
    ready_i_8_11[1] = ready_o_7_11[2];
    data_i_8_11[2] = data_o_9_11[1];
    valid_i_8_11[2] = valid_o_9_11[1];
    ready_i_8_11[2] = ready_o_9_11[1];
    data_i_8_11[0] = data_i[8][11];
    valid_i_8_11[0] = valid_i[8][11];
    ready_i_8_11[0] = ready_i[8][11];
end


/*Router 8,12*/    
merge_router #(
    .input_mask                     (input_mask_8_12),
    .output_sel                     (output_sel_8_12)
)router128(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_8_12),
    .valid_i                        (valid_i_8_12),
    .ready_o                        (ready_o_8_12),
    .data_o                         (data_o_8_12),
    .valid_o                        (valid_o_8_12),
    .ready_i                        (ready_i_8_12)
);


always@(*) begin
    data_i_8_12[3] = data_o_8_11[4];
    valid_i_8_12[3] = valid_o_8_11[4];
    ready_i_8_12[3] = ready_o_8_11[4];
    data_i_8_12[4] = data_o_8_13[3];
    valid_i_8_12[4] = valid_o_8_13[3];
    ready_i_8_12[4] = ready_o_8_13[3];
    data_i_8_12[1] = data_o_7_12[2];
    valid_i_8_12[1] = valid_o_7_12[2];
    ready_i_8_12[1] = ready_o_7_12[2];
    data_i_8_12[2] = data_o_9_12[1];
    valid_i_8_12[2] = valid_o_9_12[1];
    ready_i_8_12[2] = ready_o_9_12[1];
    data_i_8_12[0] = data_i[8][12];
    valid_i_8_12[0] = valid_i[8][12];
    ready_i_8_12[0] = ready_i[8][12];
end


/*Router 8,13*/    
merge_router #(
    .input_mask                     (input_mask_8_13),
    .output_sel                     (output_sel_8_13)
)router138(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_8_13),
    .valid_i                        (valid_i_8_13),
    .ready_o                        (ready_o_8_13),
    .data_o                         (data_o_8_13),
    .valid_o                        (valid_o_8_13),
    .ready_i                        (ready_i_8_13)
);


always@(*) begin
    data_i_8_13[3] = data_o_8_12[4];
    valid_i_8_13[3] = valid_o_8_12[4];
    ready_i_8_13[3] = ready_o_8_12[4];
    data_i_8_13[4] = data_o_8_14[3];
    valid_i_8_13[4] = valid_o_8_14[3];
    ready_i_8_13[4] = ready_o_8_14[3];
    data_i_8_13[1] = data_o_7_13[2];
    valid_i_8_13[1] = valid_o_7_13[2];
    ready_i_8_13[1] = ready_o_7_13[2];
    data_i_8_13[2] = data_o_9_13[1];
    valid_i_8_13[2] = valid_o_9_13[1];
    ready_i_8_13[2] = ready_o_9_13[1];
    data_i_8_13[0] = data_i[8][13];
    valid_i_8_13[0] = valid_i[8][13];
    ready_i_8_13[0] = ready_i[8][13];
end


/*Router 8,14*/    
merge_router #(
    .input_mask                     (input_mask_8_14),
    .output_sel                     (output_sel_8_14)
)router148(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_8_14),
    .valid_i                        (valid_i_8_14),
    .ready_o                        (ready_o_8_14),
    .data_o                         (data_o_8_14),
    .valid_o                        (valid_o_8_14),
    .ready_i                        (ready_i_8_14)
);


always@(*) begin
    data_i_8_14[3] = data_o_8_13[4];
    valid_i_8_14[3] = valid_o_8_13[4];
    ready_i_8_14[3] = ready_o_8_13[4];
    data_i_8_14[4] = data_o_8_15[3];
    valid_i_8_14[4] = valid_o_8_15[3];
    ready_i_8_14[4] = ready_o_8_15[3];
    data_i_8_14[1] = data_o_7_14[2];
    valid_i_8_14[1] = valid_o_7_14[2];
    ready_i_8_14[1] = ready_o_7_14[2];
    data_i_8_14[2] = data_o_9_14[1];
    valid_i_8_14[2] = valid_o_9_14[1];
    ready_i_8_14[2] = ready_o_9_14[1];
    data_i_8_14[0] = data_i[8][14];
    valid_i_8_14[0] = valid_i[8][14];
    ready_i_8_14[0] = ready_i[8][14];
end


/*Router 8,15*/    
merge_router #(
    .input_mask                     (input_mask_8_15),
    .output_sel                     (output_sel_8_15)
)router158(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_8_15),
    .valid_i                        (valid_i_8_15),
    .ready_o                        (ready_o_8_15),
    .data_o                         (data_o_8_15),
    .valid_o                        (valid_o_8_15),
    .ready_i                        (ready_i_8_15)
);


always@(*) begin
    data_i_8_15[3] = data_o_8_14[4];
    valid_i_8_15[3] = valid_o_8_14[4];
    ready_i_8_15[3] = ready_o_8_14[4];
    data_i_8_15[4] = data_o_8_16[3];
    valid_i_8_15[4] = valid_o_8_16[3];
    ready_i_8_15[4] = ready_o_8_16[3];
    data_i_8_15[1] = data_o_7_15[2];
    valid_i_8_15[1] = valid_o_7_15[2];
    ready_i_8_15[1] = ready_o_7_15[2];
    data_i_8_15[2] = data_o_9_15[1];
    valid_i_8_15[2] = valid_o_9_15[1];
    ready_i_8_15[2] = ready_o_9_15[1];
    data_i_8_15[0] = data_i[8][15];
    valid_i_8_15[0] = valid_i[8][15];
    ready_i_8_15[0] = ready_i[8][15];
end


/*Router 8,16*/    
merge_router #(
    .input_mask                     (input_mask_8_16),
    .output_sel                     (output_sel_8_16)
)router168(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_8_16),
    .valid_i                        (valid_i_8_16),
    .ready_o                        (ready_o_8_16),
    .data_o                         (data_o_8_16),
    .valid_o                        (valid_o_8_16),
    .ready_i                        (ready_i_8_16)
);


always@(*) begin
    data_i_8_16[3] = data_o_8_15[4];
    valid_i_8_16[3] = valid_o_8_15[4];
    ready_i_8_16[3] = ready_o_8_15[4];
    data_i_8_16[4] = data_o_8_17[3];
    valid_i_8_16[4] = valid_o_8_17[3];
    ready_i_8_16[4] = ready_o_8_17[3];
    data_i_8_16[1] = data_o_7_16[2];
    valid_i_8_16[1] = valid_o_7_16[2];
    ready_i_8_16[1] = ready_o_7_16[2];
    data_i_8_16[2] = data_o_9_16[1];
    valid_i_8_16[2] = valid_o_9_16[1];
    ready_i_8_16[2] = ready_o_9_16[1];
    data_i_8_16[0] = data_i[8][16];
    valid_i_8_16[0] = valid_i[8][16];
    ready_i_8_16[0] = ready_i[8][16];
end


/*Router 8,17*/    
merge_router #(
    .input_mask                     (input_mask_8_17),
    .output_sel                     (output_sel_8_17)
)router178(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_8_17),
    .valid_i                        (valid_i_8_17),
    .ready_o                        (ready_o_8_17),
    .data_o                         (data_o_8_17),
    .valid_o                        (valid_o_8_17),
    .ready_i                        (ready_i_8_17)
);


always@(*) begin
    data_i_8_17[3] = data_o_8_16[4];
    valid_i_8_17[3] = valid_o_8_16[4];
    ready_i_8_17[3] = ready_o_8_16[4];
    data_i_8_17[4] = data_o_8_18[3];
    valid_i_8_17[4] = valid_o_8_18[3];
    ready_i_8_17[4] = ready_o_8_18[3];
    data_i_8_17[1] = data_o_7_17[2];
    valid_i_8_17[1] = valid_o_7_17[2];
    ready_i_8_17[1] = ready_o_7_17[2];
    data_i_8_17[2] = data_o_9_17[1];
    valid_i_8_17[2] = valid_o_9_17[1];
    ready_i_8_17[2] = ready_o_9_17[1];
    data_i_8_17[0] = data_i[8][17];
    valid_i_8_17[0] = valid_i[8][17];
    ready_i_8_17[0] = ready_i[8][17];
end


/*Router 8,18*/    
merge_router #(
    .input_mask                     (input_mask_8_18),
    .output_sel                     (output_sel_8_18)
)router188(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_8_18),
    .valid_i                        (valid_i_8_18),
    .ready_o                        (ready_o_8_18),
    .data_o                         (data_o_8_18),
    .valid_o                        (valid_o_8_18),
    .ready_i                        (ready_i_8_18)
);


always@(*) begin
    data_i_8_18[3] = data_o_8_17[4];
    valid_i_8_18[3] = valid_o_8_17[4];
    ready_i_8_18[3] = ready_o_8_17[4];
    data_i_8_18[4] = data_o_8_19[3];
    valid_i_8_18[4] = valid_o_8_19[3];
    ready_i_8_18[4] = ready_o_8_19[3];
    data_i_8_18[1] = data_o_7_18[2];
    valid_i_8_18[1] = valid_o_7_18[2];
    ready_i_8_18[1] = ready_o_7_18[2];
    data_i_8_18[2] = data_o_9_18[1];
    valid_i_8_18[2] = valid_o_9_18[1];
    ready_i_8_18[2] = ready_o_9_18[1];
    data_i_8_18[0] = data_i[8][18];
    valid_i_8_18[0] = valid_i[8][18];
    ready_i_8_18[0] = ready_i[8][18];
end


/*Router 8,19*/    
merge_router #(
    .input_mask                     (input_mask_8_19),
    .output_sel                     (output_sel_8_19)
)router198(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_8_19),
    .valid_i                        (valid_i_8_19),
    .ready_o                        (ready_o_8_19),
    .data_o                         (data_o_8_19),
    .valid_o                        (valid_o_8_19),
    .ready_i                        (ready_i_8_19)
);


always@(*) begin
    data_i_8_19[3] = data_o_8_18[4];
    valid_i_8_19[3] = valid_o_8_18[4];
    ready_i_8_19[3] = ready_o_8_18[4];
    data_i_8_19[4] = data_o_8_20[3];
    valid_i_8_19[4] = valid_o_8_20[3];
    ready_i_8_19[4] = ready_o_8_20[3];
    data_i_8_19[1] = data_o_7_19[2];
    valid_i_8_19[1] = valid_o_7_19[2];
    ready_i_8_19[1] = ready_o_7_19[2];
    data_i_8_19[2] = data_o_9_19[1];
    valid_i_8_19[2] = valid_o_9_19[1];
    ready_i_8_19[2] = ready_o_9_19[1];
    data_i_8_19[0] = data_i[8][19];
    valid_i_8_19[0] = valid_i[8][19];
    ready_i_8_19[0] = ready_i[8][19];
end


/*Router 8,20*/    
merge_router #(
    .input_mask                     (input_mask_8_20),
    .output_sel                     (output_sel_8_20)
)router208(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_8_20),
    .valid_i                        (valid_i_8_20),
    .ready_o                        (ready_o_8_20),
    .data_o                         (data_o_8_20),
    .valid_o                        (valid_o_8_20),
    .ready_i                        (ready_i_8_20)
);


always@(*) begin
    data_i_8_20[3] = data_o_8_19[4];
    valid_i_8_20[3] = valid_o_8_19[4];
    ready_i_8_20[3] = ready_o_8_19[4];
    data_i_8_20[4] = data_o_8_21[3];
    valid_i_8_20[4] = valid_o_8_21[3];
    ready_i_8_20[4] = ready_o_8_21[3];
    data_i_8_20[1] = data_o_7_20[2];
    valid_i_8_20[1] = valid_o_7_20[2];
    ready_i_8_20[1] = ready_o_7_20[2];
    data_i_8_20[2] = data_o_9_20[1];
    valid_i_8_20[2] = valid_o_9_20[1];
    ready_i_8_20[2] = ready_o_9_20[1];
    data_i_8_20[0] = data_i[8][20];
    valid_i_8_20[0] = valid_i[8][20];
    ready_i_8_20[0] = ready_i[8][20];
end


/*Router 8,21*/    
merge_router #(
    .input_mask                     (input_mask_8_21),
    .output_sel                     (output_sel_8_21)
)router218(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_8_21),
    .valid_i                        (valid_i_8_21),
    .ready_o                        (ready_o_8_21),
    .data_o                         (data_o_8_21),
    .valid_o                        (valid_o_8_21),
    .ready_i                        (ready_i_8_21)
);


always@(*) begin
    data_i_8_21[3] = data_o_8_20[4];
    valid_i_8_21[3] = valid_o_8_20[4];
    ready_i_8_21[3] = ready_o_8_20[4];
    data_i_8_21[4] = data_o_8_22[3];
    valid_i_8_21[4] = valid_o_8_22[3];
    ready_i_8_21[4] = ready_o_8_22[3];
    data_i_8_21[1] = data_o_7_21[2];
    valid_i_8_21[1] = valid_o_7_21[2];
    ready_i_8_21[1] = ready_o_7_21[2];
    data_i_8_21[2] = data_o_9_21[1];
    valid_i_8_21[2] = valid_o_9_21[1];
    ready_i_8_21[2] = ready_o_9_21[1];
    data_i_8_21[0] = data_i[8][21];
    valid_i_8_21[0] = valid_i[8][21];
    ready_i_8_21[0] = ready_i[8][21];
end


/*Router 8,22*/    
merge_router #(
    .input_mask                     (input_mask_8_22),
    .output_sel                     (output_sel_8_22)
)router228(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_8_22),
    .valid_i                        (valid_i_8_22),
    .ready_o                        (ready_o_8_22),
    .data_o                         (data_o_8_22),
    .valid_o                        (valid_o_8_22),
    .ready_i                        (ready_i_8_22)
);


always@(*) begin
    data_i_8_22[3] = data_o_8_21[4];
    valid_i_8_22[3] = valid_o_8_21[4];
    ready_i_8_22[3] = ready_o_8_21[4];
    data_i_8_22[4] = data_o_8_23[3];
    valid_i_8_22[4] = valid_o_8_23[3];
    ready_i_8_22[4] = ready_o_8_23[3];
    data_i_8_22[1] = data_o_7_22[2];
    valid_i_8_22[1] = valid_o_7_22[2];
    ready_i_8_22[1] = ready_o_7_22[2];
    data_i_8_22[2] = data_o_9_22[1];
    valid_i_8_22[2] = valid_o_9_22[1];
    ready_i_8_22[2] = ready_o_9_22[1];
    data_i_8_22[0] = data_i[8][22];
    valid_i_8_22[0] = valid_i[8][22];
    ready_i_8_22[0] = ready_i[8][22];
end


/*Router 8,23*/    
merge_router #(
    .input_mask                     (input_mask_8_23),
    .output_sel                     (output_sel_8_23)
)router238(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_8_23),
    .valid_i                        (valid_i_8_23),
    .ready_o                        (ready_o_8_23),
    .data_o                         (data_o_8_23),
    .valid_o                        (valid_o_8_23),
    .ready_i                        (ready_i_8_23)
);


always@(*) begin
    data_i_8_23[3] = data_o_8_22[4];
    valid_i_8_23[3] = valid_o_8_22[4];
    ready_i_8_23[3] = ready_o_8_22[4];
    data_i_8_23[4] = data_o_8_24[3];
    valid_i_8_23[4] = valid_o_8_24[3];
    ready_i_8_23[4] = ready_o_8_24[3];
    data_i_8_23[1] = data_o_7_23[2];
    valid_i_8_23[1] = valid_o_7_23[2];
    ready_i_8_23[1] = ready_o_7_23[2];
    data_i_8_23[2] = data_o_9_23[1];
    valid_i_8_23[2] = valid_o_9_23[1];
    ready_i_8_23[2] = ready_o_9_23[1];
    data_i_8_23[0] = data_i[8][23];
    valid_i_8_23[0] = valid_i[8][23];
    ready_i_8_23[0] = ready_i[8][23];
end


/*Router 8,24*/    
merge_router #(
    .input_mask                     (input_mask_8_24),
    .output_sel                     (output_sel_8_24)
)router248(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_8_24),
    .valid_i                        (valid_i_8_24),
    .ready_o                        (ready_o_8_24),
    .data_o                         (data_o_8_24),
    .valid_o                        (valid_o_8_24),
    .ready_i                        (ready_i_8_24)
);


always@(*) begin
    data_i_8_24[3] = data_o_8_23[4];
    valid_i_8_24[3] = valid_o_8_23[4];
    ready_i_8_24[3] = ready_o_8_23[4];
    data_i_8_24[1] = data_o_7_24[2];
    valid_i_8_24[1] = valid_o_7_24[2];
    ready_i_8_24[1] = ready_o_7_24[2];
    data_i_8_24[2] = data_o_9_24[1];
    valid_i_8_24[2] = valid_o_9_24[1];
    ready_i_8_24[2] = ready_o_9_24[1];
    data_i_8_24[0] = data_i[8][24];
    valid_i_8_24[0] = valid_i[8][24];
    ready_i_8_24[0] = ready_i[8][24];
end


/*Router 9,0*/    
merge_router #(
    .input_mask                     (input_mask_9_0),
    .output_sel                     (output_sel_9_0)
)router9(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_9_0),
    .valid_i                        (valid_i_9_0),
    .ready_o                        (ready_o_9_0),
    .data_o                         (data_o_9_0),
    .valid_o                        (valid_o_9_0),
    .ready_i                        (ready_i_9_0)
);


always@(*) begin
    data_i_9_0[4] = data_o_9_1[3];
    valid_i_9_0[4] = valid_o_9_1[3];
    ready_i_9_0[4] = ready_o_9_1[3];
    data_i_9_0[1] = data_o_8_0[2];
    valid_i_9_0[1] = valid_o_8_0[2];
    ready_i_9_0[1] = ready_o_8_0[2];
    data_i_9_0[0] = data_i[9][0];
    valid_i_9_0[0] = valid_i[9][0];
    ready_i_9_0[0] = ready_i[9][0];
end


/*Router 9,1*/    
merge_router #(
    .input_mask                     (input_mask_9_1),
    .output_sel                     (output_sel_9_1)
)router19(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_9_1),
    .valid_i                        (valid_i_9_1),
    .ready_o                        (ready_o_9_1),
    .data_o                         (data_o_9_1),
    .valid_o                        (valid_o_9_1),
    .ready_i                        (ready_i_9_1)
);


always@(*) begin
    data_i_9_1[3] = data_o_9_0[4];
    valid_i_9_1[3] = valid_o_9_0[4];
    ready_i_9_1[3] = ready_o_9_0[4];
    data_i_9_1[4] = data_o_9_2[3];
    valid_i_9_1[4] = valid_o_9_2[3];
    ready_i_9_1[4] = ready_o_9_2[3];
    data_i_9_1[1] = data_o_8_1[2];
    valid_i_9_1[1] = valid_o_8_1[2];
    ready_i_9_1[1] = ready_o_8_1[2];
    data_i_9_1[0] = data_i[9][1];
    valid_i_9_1[0] = valid_i[9][1];
    ready_i_9_1[0] = ready_i[9][1];
end


/*Router 9,2*/    
merge_router #(
    .input_mask                     (input_mask_9_2),
    .output_sel                     (output_sel_9_2)
)router29(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_9_2),
    .valid_i                        (valid_i_9_2),
    .ready_o                        (ready_o_9_2),
    .data_o                         (data_o_9_2),
    .valid_o                        (valid_o_9_2),
    .ready_i                        (ready_i_9_2)
);


always@(*) begin
    data_i_9_2[3] = data_o_9_1[4];
    valid_i_9_2[3] = valid_o_9_1[4];
    ready_i_9_2[3] = ready_o_9_1[4];
    data_i_9_2[4] = data_o_9_3[3];
    valid_i_9_2[4] = valid_o_9_3[3];
    ready_i_9_2[4] = ready_o_9_3[3];
    data_i_9_2[1] = data_o_8_2[2];
    valid_i_9_2[1] = valid_o_8_2[2];
    ready_i_9_2[1] = ready_o_8_2[2];
    data_i_9_2[0] = data_i[9][2];
    valid_i_9_2[0] = valid_i[9][2];
    ready_i_9_2[0] = ready_i[9][2];
end


/*Router 9,3*/    
merge_router #(
    .input_mask                     (input_mask_9_3),
    .output_sel                     (output_sel_9_3)
)router39(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_9_3),
    .valid_i                        (valid_i_9_3),
    .ready_o                        (ready_o_9_3),
    .data_o                         (data_o_9_3),
    .valid_o                        (valid_o_9_3),
    .ready_i                        (ready_i_9_3)
);


always@(*) begin
    data_i_9_3[3] = data_o_9_2[4];
    valid_i_9_3[3] = valid_o_9_2[4];
    ready_i_9_3[3] = ready_o_9_2[4];
    data_i_9_3[4] = data_o_9_4[3];
    valid_i_9_3[4] = valid_o_9_4[3];
    ready_i_9_3[4] = ready_o_9_4[3];
    data_i_9_3[1] = data_o_8_3[2];
    valid_i_9_3[1] = valid_o_8_3[2];
    ready_i_9_3[1] = ready_o_8_3[2];
    data_i_9_3[0] = data_i[9][3];
    valid_i_9_3[0] = valid_i[9][3];
    ready_i_9_3[0] = ready_i[9][3];
end


/*Router 9,4*/    
merge_router #(
    .input_mask                     (input_mask_9_4),
    .output_sel                     (output_sel_9_4)
)router49(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_9_4),
    .valid_i                        (valid_i_9_4),
    .ready_o                        (ready_o_9_4),
    .data_o                         (data_o_9_4),
    .valid_o                        (valid_o_9_4),
    .ready_i                        (ready_i_9_4)
);


always@(*) begin
    data_i_9_4[3] = data_o_9_3[4];
    valid_i_9_4[3] = valid_o_9_3[4];
    ready_i_9_4[3] = ready_o_9_3[4];
    data_i_9_4[4] = data_o_9_5[3];
    valid_i_9_4[4] = valid_o_9_5[3];
    ready_i_9_4[4] = ready_o_9_5[3];
    data_i_9_4[1] = data_o_8_4[2];
    valid_i_9_4[1] = valid_o_8_4[2];
    ready_i_9_4[1] = ready_o_8_4[2];
    data_i_9_4[0] = data_i[9][4];
    valid_i_9_4[0] = valid_i[9][4];
    ready_i_9_4[0] = ready_i[9][4];
end


/*Router 9,5*/    
merge_router #(
    .input_mask                     (input_mask_9_5),
    .output_sel                     (output_sel_9_5)
)router59(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_9_5),
    .valid_i                        (valid_i_9_5),
    .ready_o                        (ready_o_9_5),
    .data_o                         (data_o_9_5),
    .valid_o                        (valid_o_9_5),
    .ready_i                        (ready_i_9_5)
);


always@(*) begin
    data_i_9_5[3] = data_o_9_4[4];
    valid_i_9_5[3] = valid_o_9_4[4];
    ready_i_9_5[3] = ready_o_9_4[4];
    data_i_9_5[4] = data_o_9_6[3];
    valid_i_9_5[4] = valid_o_9_6[3];
    ready_i_9_5[4] = ready_o_9_6[3];
    data_i_9_5[1] = data_o_8_5[2];
    valid_i_9_5[1] = valid_o_8_5[2];
    ready_i_9_5[1] = ready_o_8_5[2];
    data_i_9_5[0] = data_i[9][5];
    valid_i_9_5[0] = valid_i[9][5];
    ready_i_9_5[0] = ready_i[9][5];
end


/*Router 9,6*/    
merge_router #(
    .input_mask                     (input_mask_9_6),
    .output_sel                     (output_sel_9_6)
)router69(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_9_6),
    .valid_i                        (valid_i_9_6),
    .ready_o                        (ready_o_9_6),
    .data_o                         (data_o_9_6),
    .valid_o                        (valid_o_9_6),
    .ready_i                        (ready_i_9_6)
);


always@(*) begin
    data_i_9_6[3] = data_o_9_5[4];
    valid_i_9_6[3] = valid_o_9_5[4];
    ready_i_9_6[3] = ready_o_9_5[4];
    data_i_9_6[4] = data_o_9_7[3];
    valid_i_9_6[4] = valid_o_9_7[3];
    ready_i_9_6[4] = ready_o_9_7[3];
    data_i_9_6[1] = data_o_8_6[2];
    valid_i_9_6[1] = valid_o_8_6[2];
    ready_i_9_6[1] = ready_o_8_6[2];
    data_i_9_6[0] = data_i[9][6];
    valid_i_9_6[0] = valid_i[9][6];
    ready_i_9_6[0] = ready_i[9][6];
end


/*Router 9,7*/    
merge_router #(
    .input_mask                     (input_mask_9_7),
    .output_sel                     (output_sel_9_7)
)router79(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_9_7),
    .valid_i                        (valid_i_9_7),
    .ready_o                        (ready_o_9_7),
    .data_o                         (data_o_9_7),
    .valid_o                        (valid_o_9_7),
    .ready_i                        (ready_i_9_7)
);


always@(*) begin
    data_i_9_7[3] = data_o_9_6[4];
    valid_i_9_7[3] = valid_o_9_6[4];
    ready_i_9_7[3] = ready_o_9_6[4];
    data_i_9_7[4] = data_o_9_8[3];
    valid_i_9_7[4] = valid_o_9_8[3];
    ready_i_9_7[4] = ready_o_9_8[3];
    data_i_9_7[1] = data_o_8_7[2];
    valid_i_9_7[1] = valid_o_8_7[2];
    ready_i_9_7[1] = ready_o_8_7[2];
    data_i_9_7[0] = data_i[9][7];
    valid_i_9_7[0] = valid_i[9][7];
    ready_i_9_7[0] = ready_i[9][7];
end


/*Router 9,8*/    
merge_router #(
    .input_mask                     (input_mask_9_8),
    .output_sel                     (output_sel_9_8)
)router89(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_9_8),
    .valid_i                        (valid_i_9_8),
    .ready_o                        (ready_o_9_8),
    .data_o                         (data_o_9_8),
    .valid_o                        (valid_o_9_8),
    .ready_i                        (ready_i_9_8)
);


always@(*) begin
    data_i_9_8[3] = data_o_9_7[4];
    valid_i_9_8[3] = valid_o_9_7[4];
    ready_i_9_8[3] = ready_o_9_7[4];
    data_i_9_8[4] = data_o_9_9[3];
    valid_i_9_8[4] = valid_o_9_9[3];
    ready_i_9_8[4] = ready_o_9_9[3];
    data_i_9_8[1] = data_o_8_8[2];
    valid_i_9_8[1] = valid_o_8_8[2];
    ready_i_9_8[1] = ready_o_8_8[2];
    data_i_9_8[0] = data_i[9][8];
    valid_i_9_8[0] = valid_i[9][8];
    ready_i_9_8[0] = ready_i[9][8];
end


/*Router 9,9*/    
merge_router #(
    .input_mask                     (input_mask_9_9),
    .output_sel                     (output_sel_9_9)
)router99(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_9_9),
    .valid_i                        (valid_i_9_9),
    .ready_o                        (ready_o_9_9),
    .data_o                         (data_o_9_9),
    .valid_o                        (valid_o_9_9),
    .ready_i                        (ready_i_9_9)
);


always@(*) begin
    data_i_9_9[3] = data_o_9_8[4];
    valid_i_9_9[3] = valid_o_9_8[4];
    ready_i_9_9[3] = ready_o_9_8[4];
    data_i_9_9[4] = data_o_9_10[3];
    valid_i_9_9[4] = valid_o_9_10[3];
    ready_i_9_9[4] = ready_o_9_10[3];
    data_i_9_9[1] = data_o_8_9[2];
    valid_i_9_9[1] = valid_o_8_9[2];
    ready_i_9_9[1] = ready_o_8_9[2];
    data_i_9_9[0] = data_i[9][9];
    valid_i_9_9[0] = valid_i[9][9];
    ready_i_9_9[0] = ready_i[9][9];
end


/*Router 9,10*/    
merge_router #(
    .input_mask                     (input_mask_9_10),
    .output_sel                     (output_sel_9_10)
)router109(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_9_10),
    .valid_i                        (valid_i_9_10),
    .ready_o                        (ready_o_9_10),
    .data_o                         (data_o_9_10),
    .valid_o                        (valid_o_9_10),
    .ready_i                        (ready_i_9_10)
);


always@(*) begin
    data_i_9_10[3] = data_o_9_9[4];
    valid_i_9_10[3] = valid_o_9_9[4];
    ready_i_9_10[3] = ready_o_9_9[4];
    data_i_9_10[4] = data_o_9_11[3];
    valid_i_9_10[4] = valid_o_9_11[3];
    ready_i_9_10[4] = ready_o_9_11[3];
    data_i_9_10[1] = data_o_8_10[2];
    valid_i_9_10[1] = valid_o_8_10[2];
    ready_i_9_10[1] = ready_o_8_10[2];
    data_i_9_10[0] = data_i[9][10];
    valid_i_9_10[0] = valid_i[9][10];
    ready_i_9_10[0] = ready_i[9][10];
end


/*Router 9,11*/    
merge_router #(
    .input_mask                     (input_mask_9_11),
    .output_sel                     (output_sel_9_11)
)router119(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_9_11),
    .valid_i                        (valid_i_9_11),
    .ready_o                        (ready_o_9_11),
    .data_o                         (data_o_9_11),
    .valid_o                        (valid_o_9_11),
    .ready_i                        (ready_i_9_11)
);


always@(*) begin
    data_i_9_11[3] = data_o_9_10[4];
    valid_i_9_11[3] = valid_o_9_10[4];
    ready_i_9_11[3] = ready_o_9_10[4];
    data_i_9_11[4] = data_o_9_12[3];
    valid_i_9_11[4] = valid_o_9_12[3];
    ready_i_9_11[4] = ready_o_9_12[3];
    data_i_9_11[1] = data_o_8_11[2];
    valid_i_9_11[1] = valid_o_8_11[2];
    ready_i_9_11[1] = ready_o_8_11[2];
    data_i_9_11[0] = data_i[9][11];
    valid_i_9_11[0] = valid_i[9][11];
    ready_i_9_11[0] = ready_i[9][11];
end


/*Router 9,12*/    
merge_router #(
    .input_mask                     (input_mask_9_12),
    .output_sel                     (output_sel_9_12)
)router129(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_9_12),
    .valid_i                        (valid_i_9_12),
    .ready_o                        (ready_o_9_12),
    .data_o                         (data_o_9_12),
    .valid_o                        (valid_o_9_12),
    .ready_i                        (ready_i_9_12)
);


always@(*) begin
    data_i_9_12[3] = data_o_9_11[4];
    valid_i_9_12[3] = valid_o_9_11[4];
    ready_i_9_12[3] = ready_o_9_11[4];
    data_i_9_12[4] = data_o_9_13[3];
    valid_i_9_12[4] = valid_o_9_13[3];
    ready_i_9_12[4] = ready_o_9_13[3];
    data_i_9_12[1] = data_o_8_12[2];
    valid_i_9_12[1] = valid_o_8_12[2];
    ready_i_9_12[1] = ready_o_8_12[2];
    data_i_9_12[0] = data_i[9][12];
    valid_i_9_12[0] = valid_i[9][12];
    ready_i_9_12[0] = ready_i[9][12];
end


/*Router 9,13*/    
merge_router #(
    .input_mask                     (input_mask_9_13),
    .output_sel                     (output_sel_9_13)
)router139(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_9_13),
    .valid_i                        (valid_i_9_13),
    .ready_o                        (ready_o_9_13),
    .data_o                         (data_o_9_13),
    .valid_o                        (valid_o_9_13),
    .ready_i                        (ready_i_9_13)
);


always@(*) begin
    data_i_9_13[3] = data_o_9_12[4];
    valid_i_9_13[3] = valid_o_9_12[4];
    ready_i_9_13[3] = ready_o_9_12[4];
    data_i_9_13[4] = data_o_9_14[3];
    valid_i_9_13[4] = valid_o_9_14[3];
    ready_i_9_13[4] = ready_o_9_14[3];
    data_i_9_13[1] = data_o_8_13[2];
    valid_i_9_13[1] = valid_o_8_13[2];
    ready_i_9_13[1] = ready_o_8_13[2];
    data_i_9_13[0] = data_i[9][13];
    valid_i_9_13[0] = valid_i[9][13];
    ready_i_9_13[0] = ready_i[9][13];
end


/*Router 9,14*/    
merge_router #(
    .input_mask                     (input_mask_9_14),
    .output_sel                     (output_sel_9_14)
)router149(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_9_14),
    .valid_i                        (valid_i_9_14),
    .ready_o                        (ready_o_9_14),
    .data_o                         (data_o_9_14),
    .valid_o                        (valid_o_9_14),
    .ready_i                        (ready_i_9_14)
);


always@(*) begin
    data_i_9_14[3] = data_o_9_13[4];
    valid_i_9_14[3] = valid_o_9_13[4];
    ready_i_9_14[3] = ready_o_9_13[4];
    data_i_9_14[4] = data_o_9_15[3];
    valid_i_9_14[4] = valid_o_9_15[3];
    ready_i_9_14[4] = ready_o_9_15[3];
    data_i_9_14[1] = data_o_8_14[2];
    valid_i_9_14[1] = valid_o_8_14[2];
    ready_i_9_14[1] = ready_o_8_14[2];
    data_i_9_14[0] = data_i[9][14];
    valid_i_9_14[0] = valid_i[9][14];
    ready_i_9_14[0] = ready_i[9][14];
end


/*Router 9,15*/    
merge_router #(
    .input_mask                     (input_mask_9_15),
    .output_sel                     (output_sel_9_15)
)router159(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_9_15),
    .valid_i                        (valid_i_9_15),
    .ready_o                        (ready_o_9_15),
    .data_o                         (data_o_9_15),
    .valid_o                        (valid_o_9_15),
    .ready_i                        (ready_i_9_15)
);


always@(*) begin
    data_i_9_15[3] = data_o_9_14[4];
    valid_i_9_15[3] = valid_o_9_14[4];
    ready_i_9_15[3] = ready_o_9_14[4];
    data_i_9_15[4] = data_o_9_16[3];
    valid_i_9_15[4] = valid_o_9_16[3];
    ready_i_9_15[4] = ready_o_9_16[3];
    data_i_9_15[1] = data_o_8_15[2];
    valid_i_9_15[1] = valid_o_8_15[2];
    ready_i_9_15[1] = ready_o_8_15[2];
    data_i_9_15[0] = data_i[9][15];
    valid_i_9_15[0] = valid_i[9][15];
    ready_i_9_15[0] = ready_i[9][15];
end


/*Router 9,16*/    
merge_router #(
    .input_mask                     (input_mask_9_16),
    .output_sel                     (output_sel_9_16)
)router169(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_9_16),
    .valid_i                        (valid_i_9_16),
    .ready_o                        (ready_o_9_16),
    .data_o                         (data_o_9_16),
    .valid_o                        (valid_o_9_16),
    .ready_i                        (ready_i_9_16)
);


always@(*) begin
    data_i_9_16[3] = data_o_9_15[4];
    valid_i_9_16[3] = valid_o_9_15[4];
    ready_i_9_16[3] = ready_o_9_15[4];
    data_i_9_16[4] = data_o_9_17[3];
    valid_i_9_16[4] = valid_o_9_17[3];
    ready_i_9_16[4] = ready_o_9_17[3];
    data_i_9_16[1] = data_o_8_16[2];
    valid_i_9_16[1] = valid_o_8_16[2];
    ready_i_9_16[1] = ready_o_8_16[2];
    data_i_9_16[0] = data_i[9][16];
    valid_i_9_16[0] = valid_i[9][16];
    ready_i_9_16[0] = ready_i[9][16];
end


/*Router 9,17*/    
merge_router #(
    .input_mask                     (input_mask_9_17),
    .output_sel                     (output_sel_9_17)
)router179(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_9_17),
    .valid_i                        (valid_i_9_17),
    .ready_o                        (ready_o_9_17),
    .data_o                         (data_o_9_17),
    .valid_o                        (valid_o_9_17),
    .ready_i                        (ready_i_9_17)
);


always@(*) begin
    data_i_9_17[3] = data_o_9_16[4];
    valid_i_9_17[3] = valid_o_9_16[4];
    ready_i_9_17[3] = ready_o_9_16[4];
    data_i_9_17[4] = data_o_9_18[3];
    valid_i_9_17[4] = valid_o_9_18[3];
    ready_i_9_17[4] = ready_o_9_18[3];
    data_i_9_17[1] = data_o_8_17[2];
    valid_i_9_17[1] = valid_o_8_17[2];
    ready_i_9_17[1] = ready_o_8_17[2];
    data_i_9_17[0] = data_i[9][17];
    valid_i_9_17[0] = valid_i[9][17];
    ready_i_9_17[0] = ready_i[9][17];
end


/*Router 9,18*/    
merge_router #(
    .input_mask                     (input_mask_9_18),
    .output_sel                     (output_sel_9_18)
)router189(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_9_18),
    .valid_i                        (valid_i_9_18),
    .ready_o                        (ready_o_9_18),
    .data_o                         (data_o_9_18),
    .valid_o                        (valid_o_9_18),
    .ready_i                        (ready_i_9_18)
);


always@(*) begin
    data_i_9_18[3] = data_o_9_17[4];
    valid_i_9_18[3] = valid_o_9_17[4];
    ready_i_9_18[3] = ready_o_9_17[4];
    data_i_9_18[4] = data_o_9_19[3];
    valid_i_9_18[4] = valid_o_9_19[3];
    ready_i_9_18[4] = ready_o_9_19[3];
    data_i_9_18[1] = data_o_8_18[2];
    valid_i_9_18[1] = valid_o_8_18[2];
    ready_i_9_18[1] = ready_o_8_18[2];
    data_i_9_18[0] = data_i[9][18];
    valid_i_9_18[0] = valid_i[9][18];
    ready_i_9_18[0] = ready_i[9][18];
end


/*Router 9,19*/    
merge_router #(
    .input_mask                     (input_mask_9_19),
    .output_sel                     (output_sel_9_19)
)router199(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_9_19),
    .valid_i                        (valid_i_9_19),
    .ready_o                        (ready_o_9_19),
    .data_o                         (data_o_9_19),
    .valid_o                        (valid_o_9_19),
    .ready_i                        (ready_i_9_19)
);


always@(*) begin
    data_i_9_19[3] = data_o_9_18[4];
    valid_i_9_19[3] = valid_o_9_18[4];
    ready_i_9_19[3] = ready_o_9_18[4];
    data_i_9_19[4] = data_o_9_20[3];
    valid_i_9_19[4] = valid_o_9_20[3];
    ready_i_9_19[4] = ready_o_9_20[3];
    data_i_9_19[1] = data_o_8_19[2];
    valid_i_9_19[1] = valid_o_8_19[2];
    ready_i_9_19[1] = ready_o_8_19[2];
    data_i_9_19[0] = data_i[9][19];
    valid_i_9_19[0] = valid_i[9][19];
    ready_i_9_19[0] = ready_i[9][19];
end


/*Router 9,20*/    
merge_router #(
    .input_mask                     (input_mask_9_20),
    .output_sel                     (output_sel_9_20)
)router209(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_9_20),
    .valid_i                        (valid_i_9_20),
    .ready_o                        (ready_o_9_20),
    .data_o                         (data_o_9_20),
    .valid_o                        (valid_o_9_20),
    .ready_i                        (ready_i_9_20)
);


always@(*) begin
    data_i_9_20[3] = data_o_9_19[4];
    valid_i_9_20[3] = valid_o_9_19[4];
    ready_i_9_20[3] = ready_o_9_19[4];
    data_i_9_20[4] = data_o_9_21[3];
    valid_i_9_20[4] = valid_o_9_21[3];
    ready_i_9_20[4] = ready_o_9_21[3];
    data_i_9_20[1] = data_o_8_20[2];
    valid_i_9_20[1] = valid_o_8_20[2];
    ready_i_9_20[1] = ready_o_8_20[2];
    data_i_9_20[0] = data_i[9][20];
    valid_i_9_20[0] = valid_i[9][20];
    ready_i_9_20[0] = ready_i[9][20];
end


/*Router 9,21*/    
merge_router #(
    .input_mask                     (input_mask_9_21),
    .output_sel                     (output_sel_9_21)
)router219(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_9_21),
    .valid_i                        (valid_i_9_21),
    .ready_o                        (ready_o_9_21),
    .data_o                         (data_o_9_21),
    .valid_o                        (valid_o_9_21),
    .ready_i                        (ready_i_9_21)
);


always@(*) begin
    data_i_9_21[3] = data_o_9_20[4];
    valid_i_9_21[3] = valid_o_9_20[4];
    ready_i_9_21[3] = ready_o_9_20[4];
    data_i_9_21[4] = data_o_9_22[3];
    valid_i_9_21[4] = valid_o_9_22[3];
    ready_i_9_21[4] = ready_o_9_22[3];
    data_i_9_21[1] = data_o_8_21[2];
    valid_i_9_21[1] = valid_o_8_21[2];
    ready_i_9_21[1] = ready_o_8_21[2];
    data_i_9_21[0] = data_i[9][21];
    valid_i_9_21[0] = valid_i[9][21];
    ready_i_9_21[0] = ready_i[9][21];
end


/*Router 9,22*/    
merge_router #(
    .input_mask                     (input_mask_9_22),
    .output_sel                     (output_sel_9_22)
)router229(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_9_22),
    .valid_i                        (valid_i_9_22),
    .ready_o                        (ready_o_9_22),
    .data_o                         (data_o_9_22),
    .valid_o                        (valid_o_9_22),
    .ready_i                        (ready_i_9_22)
);


always@(*) begin
    data_i_9_22[3] = data_o_9_21[4];
    valid_i_9_22[3] = valid_o_9_21[4];
    ready_i_9_22[3] = ready_o_9_21[4];
    data_i_9_22[4] = data_o_9_23[3];
    valid_i_9_22[4] = valid_o_9_23[3];
    ready_i_9_22[4] = ready_o_9_23[3];
    data_i_9_22[1] = data_o_8_22[2];
    valid_i_9_22[1] = valid_o_8_22[2];
    ready_i_9_22[1] = ready_o_8_22[2];
    data_i_9_22[0] = data_i[9][22];
    valid_i_9_22[0] = valid_i[9][22];
    ready_i_9_22[0] = ready_i[9][22];
end


/*Router 9,23*/    
merge_router #(
    .input_mask                     (input_mask_9_23),
    .output_sel                     (output_sel_9_23)
)router239(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_9_23),
    .valid_i                        (valid_i_9_23),
    .ready_o                        (ready_o_9_23),
    .data_o                         (data_o_9_23),
    .valid_o                        (valid_o_9_23),
    .ready_i                        (ready_i_9_23)
);


always@(*) begin
    data_i_9_23[3] = data_o_9_22[4];
    valid_i_9_23[3] = valid_o_9_22[4];
    ready_i_9_23[3] = ready_o_9_22[4];
    data_i_9_23[4] = data_o_9_24[3];
    valid_i_9_23[4] = valid_o_9_24[3];
    ready_i_9_23[4] = ready_o_9_24[3];
    data_i_9_23[1] = data_o_8_23[2];
    valid_i_9_23[1] = valid_o_8_23[2];
    ready_i_9_23[1] = ready_o_8_23[2];
    data_i_9_23[0] = data_i[9][23];
    valid_i_9_23[0] = valid_i[9][23];
    ready_i_9_23[0] = ready_i[9][23];
end


/*Router 9,24*/    
merge_router #(
    .input_mask                     (input_mask_9_24),
    .output_sel                     (output_sel_9_24)
)router249(
    .clk                            (clk),
    .rstn                           (rstn),
    .data_i                         (data_i_9_24),
    .valid_i                        (valid_i_9_24),
    .ready_o                        (ready_o_9_24),
    .data_o                         (data_o_9_24),
    .valid_o                        (valid_o_9_24),
    .ready_i                        (ready_i_9_24)
);


always@(*) begin
    data_i_9_24[3] = data_o_9_23[4];
    valid_i_9_24[3] = valid_o_9_23[4];
    ready_i_9_24[3] = ready_o_9_23[4];
    data_i_9_24[1] = data_o_8_24[2];
    valid_i_9_24[1] = valid_o_8_24[2];
    ready_i_9_24[1] = ready_o_8_24[2];
    data_i_9_24[0] = data_i[9][24];
    valid_i_9_24[0] = valid_i[9][24];
    ready_i_9_24[0] = ready_i[9][24];
end


endmodule
