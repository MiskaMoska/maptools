localparam isUBM_list_0_0[`CN] = '{1,1,1,1,1};
localparam isUBM_list_1_0[`CN] = '{1,1,1,1,1};
localparam isUBM_list_2_0[`CN] = '{1,1,1,1,1};
localparam isUBM_list_0_1[`CN] = '{1,1,1,1,1};
localparam isUBM_list_1_1[`CN] = '{1,1,1,1,1};
localparam isUBM_list_2_1[`CN] = '{1,1,1,1,1};
localparam isUBM_list_0_2[`CN] = '{1,1,1,1,1};
localparam isUBM_list_1_2[`CN] = '{1,1,1,1,1};
localparam isUBM_list_2_2[`CN] = '{1,1,1,1,1};

localparam isFC_list_0_0[`CN] = '{0,0,0,0,0};
localparam isFC_list_1_0[`CN] = '{1,0,0,0,0};
localparam isFC_list_2_0[`CN] = '{1,0,0,0,0};
localparam isFC_list_0_1[`CN] = '{0,0,0,0,0};
localparam isFC_list_1_1[`CN] = '{0,0,0,0,0};
localparam isFC_list_2_1[`CN] = '{0,0,0,0,0};
localparam isFC_list_0_2[`CN] = '{0,0,0,0,0};
localparam isFC_list_1_2[`CN] = '{0,0,0,0,0};
localparam isFC_list_2_2[`CN] = '{0,0,0,0,0};

localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_0_0[`CN] = '{9'b0,9'b0,9'b0,9'b0,9'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_1_0[`CN] = '{9'b100010100,9'b0,9'b0,9'b0,9'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_2_0[`CN] = '{9'b011101011,9'b0,9'b0,9'b0,9'b0}; //note the reverse index
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_0_1[`CN] = '{9'b0,9'b0,9'b0,9'b0,9'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_1_1[`CN] = '{9'b0,9'b0,9'b0,9'b0,9'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_2_1[`CN] = '{9'b0,9'b0,9'b0,9'b0,9'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_0_2[`CN] = '{9'b0,9'b0,9'b0,9'b0,9'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_1_2[`CN] = '{9'b0,9'b0,9'b0,9'b0,9'b0};
localparam [`NOC_WIDTH*`NOC_HEIGHT-1:0] FCdn_list_2_2[`CN] = '{9'b0,9'b0,9'b0,9'b0,9'b0};

localparam int FCpl_list_0_0[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_1_0[`CN] = '{16,0,0,0,0};
localparam int FCpl_list_2_0[`CN] = '{16,0,0,0,0};
localparam int FCpl_list_0_1[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_1_1[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_2_1[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_0_2[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_1_2[`CN] = '{0,0,0,0,0};
localparam int FCpl_list_2_2[`CN] = '{0,0,0,0,0};

localparam string rt_file_list_0_0[`CN] = '{"/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_0_0_0","/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_0_0_1","/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_0_0_2","/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_0_0_3","/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_0_0_4"};
localparam string rt_file_list_1_0[`CN] = '{"/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_1_0_0","/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_1_0_1","/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_1_0_2","/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_1_0_3","/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_1_0_4"};
localparam string rt_file_list_2_0[`CN] = '{"/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_2_0_0","/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_2_0_1","/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_2_0_2","/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_2_0_3","/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_2_0_4"};
localparam string rt_file_list_0_1[`CN] = '{"/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_0_1_0","/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_0_1_1","/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_0_1_2","/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_0_1_3","/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_0_1_4"};
localparam string rt_file_list_1_1[`CN] = '{"/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_1_1_0","/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_1_1_1","/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_1_1_2","/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_1_1_3","/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_1_1_4"};
localparam string rt_file_list_2_1[`CN] = '{"/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_2_1_0","/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_2_1_1","/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_2_1_2","/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_2_1_3","/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_2_1_4"};
localparam string rt_file_list_0_2[`CN] = '{"/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_0_2_0","/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_0_2_1","/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_0_2_2","/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_0_2_3","/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_0_2_4"};
localparam string rt_file_list_1_2[`CN] = '{"/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_1_2_0","/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_1_2_1","/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_1_2_2","/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_1_2_3","/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_1_2_4"};
localparam string rt_file_list_2_2[`CN] = '{"/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_2_2_0","/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_2_2_1","/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_2_2_2","/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_2_2_3","/mnt/c/git/NVCIM-COMM/behavior_model/test_dual_multicast/config/cast_rt_2_2_4"};
