localparam input_mask_0_0 = 5'b00000;
localparam output_sel_0_0 = 5'b00001;
localparam input_mask_0_1 = 5'b00001;
localparam output_sel_0_1 = 5'b10000;
localparam input_mask_0_2 = 5'b01001;
localparam output_sel_0_2 = 5'b00100;
localparam input_mask_0_3 = 5'b00101;
localparam output_sel_0_3 = 5'b10000;
localparam input_mask_0_4 = 5'b01000;
localparam output_sel_0_4 = 5'b00001;
localparam input_mask_0_5 = 5'b00001;
localparam output_sel_0_5 = 5'b10000;
localparam input_mask_0_6 = 5'b01100;
localparam output_sel_0_6 = 5'b00001;
localparam input_mask_0_7 = 5'b00000;
localparam output_sel_0_7 = 5'b00001;
localparam input_mask_1_0 = 5'b00000;
localparam output_sel_1_0 = 5'b00001;
localparam input_mask_1_1 = 5'b00100;
localparam output_sel_1_1 = 5'b00001;
localparam input_mask_1_2 = 5'b00110;
localparam output_sel_1_2 = 5'b00001;
localparam input_mask_1_3 = 5'b00101;
localparam output_sel_1_3 = 5'b00010;
localparam input_mask_1_4 = 5'b00001;
localparam output_sel_1_4 = 5'b00100;
localparam input_mask_1_5 = 5'b00001;
localparam output_sel_1_5 = 5'b10000;
localparam input_mask_1_6 = 5'b01001;
localparam output_sel_1_6 = 5'b00010;
localparam input_mask_1_7 = 5'b00000;
localparam output_sel_1_7 = 5'b00001;
localparam input_mask_2_0 = 5'b00000;
localparam output_sel_2_0 = 5'b00001;
localparam input_mask_2_1 = 5'b00001;
localparam output_sel_2_1 = 5'b00010;
localparam input_mask_2_2 = 5'b00001;
localparam output_sel_2_2 = 5'b00010;
localparam input_mask_2_3 = 5'b00001;
localparam output_sel_2_3 = 5'b00010;
localparam input_mask_2_4 = 5'b00011;
localparam output_sel_2_4 = 5'b00100;
localparam input_mask_2_5 = 5'b00101;
localparam output_sel_2_5 = 5'b10000;
localparam input_mask_2_6 = 5'b01000;
localparam output_sel_2_6 = 5'b00001;
localparam input_mask_2_7 = 5'b00000;
localparam output_sel_2_7 = 5'b00001;
localparam input_mask_3_0 = 5'b00000;
localparam output_sel_3_0 = 5'b00001;
localparam input_mask_3_1 = 5'b00100;
localparam output_sel_3_1 = 5'b00001;
localparam input_mask_3_2 = 5'b00001;
localparam output_sel_3_2 = 5'b00100;
localparam input_mask_3_3 = 5'b00100;
localparam output_sel_3_3 = 5'b00001;
localparam input_mask_3_4 = 5'b00011;
localparam output_sel_3_4 = 5'b00100;
localparam input_mask_3_5 = 5'b00101;
localparam output_sel_3_5 = 5'b00010;
localparam input_mask_3_6 = 5'b00001;
localparam output_sel_3_6 = 5'b10000;
localparam input_mask_3_7 = 5'b01100;
localparam output_sel_3_7 = 5'b00001;
localparam input_mask_4_0 = 5'b00000;
localparam output_sel_4_0 = 5'b00001;
localparam input_mask_4_1 = 5'b00001;
localparam output_sel_4_1 = 5'b00010;
localparam input_mask_4_2 = 5'b00110;
localparam output_sel_4_2 = 5'b00001;
localparam input_mask_4_3 = 5'b00101;
localparam output_sel_4_3 = 5'b00010;
localparam input_mask_4_4 = 5'b00010;
localparam output_sel_4_4 = 5'b00001;
localparam input_mask_4_5 = 5'b00001;
localparam output_sel_4_5 = 5'b00010;
localparam input_mask_4_6 = 5'b00001;
localparam output_sel_4_6 = 5'b10000;
localparam input_mask_4_7 = 5'b01001;
localparam output_sel_4_7 = 5'b00010;
localparam input_mask_5_0 = 5'b00001;
localparam output_sel_5_0 = 5'b00100;
localparam input_mask_5_1 = 5'b00100;
localparam output_sel_5_1 = 5'b00001;
localparam input_mask_5_2 = 5'b00101;
localparam output_sel_5_2 = 5'b00010;
localparam input_mask_5_3 = 5'b00101;
localparam output_sel_5_3 = 5'b00010;
localparam input_mask_5_4 = 5'b00001;
localparam output_sel_5_4 = 5'b10000;
localparam input_mask_5_5 = 5'b01100;
localparam output_sel_5_5 = 5'b00001;
localparam input_mask_5_6 = 5'b00001;
localparam output_sel_5_6 = 5'b10000;
localparam input_mask_5_7 = 5'b01100;
localparam output_sel_5_7 = 5'b00001;
localparam input_mask_6_0 = 5'b00010;
localparam output_sel_6_0 = 5'b00001;
localparam input_mask_6_1 = 5'b00001;
localparam output_sel_6_1 = 5'b00010;
localparam input_mask_6_2 = 5'b00001;
localparam output_sel_6_2 = 5'b00010;
localparam input_mask_6_3 = 5'b00001;
localparam output_sel_6_3 = 5'b00010;
localparam input_mask_6_4 = 5'b00001;
localparam output_sel_6_4 = 5'b10000;
localparam input_mask_6_5 = 5'b01001;
localparam output_sel_6_5 = 5'b00010;
localparam input_mask_6_6 = 5'b00001;
localparam output_sel_6_6 = 5'b10000;
localparam input_mask_6_7 = 5'b01001;
localparam output_sel_6_7 = 5'b00010;