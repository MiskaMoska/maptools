localparam isPooler_0_0 = 0;
localparam isCaster_0_0 = 1;
localparam stream_id_0_0 = 1;
localparam isPooler_0_1 = 0;
localparam isCaster_0_1 = 0;
localparam stream_id_0_1 = 0;
localparam isPooler_0_2 = 0;
localparam isCaster_0_2 = 1;
localparam stream_id_0_2 = 8;
localparam isPooler_0_3 = 0;
localparam isCaster_0_3 = 0;
localparam stream_id_0_3 = 0;
localparam isPooler_0_4 = 0;
localparam isCaster_0_4 = 1;
localparam stream_id_0_4 = 11;
localparam isPooler_0_5 = 0;
localparam isCaster_0_5 = 0;
localparam stream_id_0_5 = 0;
localparam isPooler_0_6 = 0;
localparam isCaster_0_6 = 0;
localparam stream_id_0_6 = 0;
localparam isPooler_0_7 = 0;
localparam isCaster_0_7 = 0;
localparam stream_id_0_7 = 0;
localparam isPooler_0_8 = 0;
localparam isCaster_0_8 = 1;
localparam stream_id_0_8 = 16;
localparam isPooler_0_9 = 0;
localparam isCaster_0_9 = 0;
localparam stream_id_0_9 = 0;
localparam isPooler_0_10 = 0;
localparam isCaster_0_10 = 0;
localparam stream_id_0_10 = 0;
localparam isPooler_1_0 = 0;
localparam isCaster_1_0 = 1;
localparam stream_id_1_0 = 2;
localparam isPooler_1_1 = 0;
localparam isCaster_1_1 = 1;
localparam stream_id_1_1 = 7;
localparam isPooler_1_2 = 0;
localparam isCaster_1_2 = 0;
localparam stream_id_1_2 = 0;
localparam isPooler_1_3 = 0;
localparam isCaster_1_3 = 0;
localparam stream_id_1_3 = 0;
localparam isPooler_1_4 = 0;
localparam isCaster_1_4 = 0;
localparam stream_id_1_4 = 0;
localparam isPooler_1_5 = 0;
localparam isCaster_1_5 = 1;
localparam stream_id_1_5 = 13;
localparam isPooler_1_6 = 0;
localparam isCaster_1_6 = 1;
localparam stream_id_1_6 = 14;
localparam isPooler_1_7 = 0;
localparam isCaster_1_7 = 0;
localparam stream_id_1_7 = 0;
localparam isPooler_1_8 = 0;
localparam isCaster_1_8 = 0;
localparam stream_id_1_8 = 0;
localparam isPooler_1_9 = 0;
localparam isCaster_1_9 = 0;
localparam stream_id_1_9 = 0;
localparam isPooler_1_10 = 0;
localparam isCaster_1_10 = 1;
localparam stream_id_1_10 = 1022;
localparam isPooler_2_0 = 1;
localparam isCaster_2_0 = 1;
localparam stream_id_2_0 = 3;
localparam isPooler_2_1 = 0;
localparam isCaster_2_1 = 0;
localparam stream_id_2_1 = 0;
localparam isPooler_2_2 = 0;
localparam isCaster_2_2 = 1;
localparam stream_id_2_2 = 9;
localparam isPooler_2_3 = 0;
localparam isCaster_2_3 = 0;
localparam stream_id_2_3 = 0;
localparam isPooler_2_4 = 0;
localparam isCaster_2_4 = 1;
localparam stream_id_2_4 = 12;
localparam isPooler_2_5 = 0;
localparam isCaster_2_5 = 0;
localparam stream_id_2_5 = 0;
localparam isPooler_2_6 = 0;
localparam isCaster_2_6 = 0;
localparam stream_id_2_6 = 0;
localparam isPooler_2_7 = 0;
localparam isCaster_2_7 = 0;
localparam stream_id_2_7 = 0;
localparam isPooler_2_8 = 0;
localparam isCaster_2_8 = 0;
localparam stream_id_2_8 = 0;
localparam isPooler_2_9 = 0;
localparam isCaster_2_9 = 0;
localparam stream_id_2_9 = 0;
localparam isPooler_2_10 = 0;
localparam isCaster_2_10 = 0;
localparam stream_id_2_10 = 0;
localparam isPooler_3_0 = 0;
localparam isCaster_3_0 = 1;
localparam stream_id_3_0 = 4;
localparam isPooler_3_1 = 0;
localparam isCaster_3_1 = 1;
localparam stream_id_3_1 = 6;
localparam isPooler_3_2 = 0;
localparam isCaster_3_2 = 0;
localparam stream_id_3_2 = 0;
localparam isPooler_3_3 = 0;
localparam isCaster_3_3 = 0;
localparam stream_id_3_3 = 0;
localparam isPooler_3_4 = 0;
localparam isCaster_3_4 = 0;
localparam stream_id_3_4 = 0;
localparam isPooler_3_5 = 0;
localparam isCaster_3_5 = 0;
localparam stream_id_3_5 = 0;
localparam isPooler_3_6 = 0;
localparam isCaster_3_6 = 0;
localparam stream_id_3_6 = 0;
localparam isPooler_3_7 = 0;
localparam isCaster_3_7 = 0;
localparam stream_id_3_7 = 0;
localparam isPooler_3_8 = 0;
localparam isCaster_3_8 = 1;
localparam stream_id_3_8 = 17;
localparam isPooler_3_9 = 0;
localparam isCaster_3_9 = 1;
localparam stream_id_3_9 = 1022;
localparam isPooler_3_10 = 0;
localparam isCaster_3_10 = 0;
localparam stream_id_3_10 = 0;
localparam isPooler_4_0 = 0;
localparam isCaster_4_0 = 1;
localparam stream_id_4_0 = 5;
localparam isPooler_4_1 = 0;
localparam isCaster_4_1 = 0;
localparam stream_id_4_1 = 0;
localparam isPooler_4_2 = 0;
localparam isCaster_4_2 = 0;
localparam stream_id_4_2 = 0;
localparam isPooler_4_3 = 0;
localparam isCaster_4_3 = 1;
localparam stream_id_4_3 = 10;
localparam isPooler_4_4 = 0;
localparam isCaster_4_4 = 0;
localparam stream_id_4_4 = 0;
localparam isPooler_4_5 = 0;
localparam isCaster_4_5 = 0;
localparam stream_id_4_5 = 0;
localparam isPooler_4_6 = 0;
localparam isCaster_4_6 = 0;
localparam stream_id_4_6 = 0;
localparam isPooler_4_7 = 0;
localparam isCaster_4_7 = 1;
localparam stream_id_4_7 = 15;
localparam isPooler_4_8 = 0;
localparam isCaster_4_8 = 0;
localparam stream_id_4_8 = 0;
localparam isPooler_4_9 = 0;
localparam isCaster_4_9 = 0;
localparam stream_id_4_9 = 0;
localparam isPooler_4_10 = 0;
localparam isCaster_4_10 = 0;
localparam stream_id_4_10 = 0;

