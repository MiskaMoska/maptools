
`ifndef __NETWORK_CONFIG_SVH_
`define __NETWORK_CONFIG_SVH_
    
localparam cast_out_0_0 = 1;
localparam merge_out_0_0 = 0;
localparam gather_out_0_0 = 1;
localparam merge_in_0_0 = 0;
localparam gather_in_0_0 = 0;
localparam cast_sid_0_0 = 1;
localparam gather_sid_0_0 = 1;

localparam cast_out_0_1 = 1;
localparam merge_out_0_1 = 0;
localparam gather_out_0_1 = 0;
localparam merge_in_0_1 = 0;
localparam gather_in_0_1 = 1;
localparam cast_sid_0_1 = 9;
localparam gather_sid_0_1 = 0;

localparam cast_out_0_2 = 1;
localparam merge_out_0_2 = 0;
localparam gather_out_0_2 = 0;
localparam merge_in_0_2 = 0;
localparam gather_in_0_2 = 0;
localparam cast_sid_0_2 = 10;
localparam gather_sid_0_2 = 0;

localparam cast_out_0_3 = 1;
localparam merge_out_0_3 = 0;
localparam gather_out_0_3 = 0;
localparam merge_in_0_3 = 1;
localparam gather_in_0_3 = 0;
localparam cast_sid_0_3 = 14;
localparam gather_sid_0_3 = 0;

localparam cast_out_0_4 = 0;
localparam merge_out_0_4 = 1;
localparam gather_out_0_4 = 0;
localparam merge_in_0_4 = 0;
localparam gather_in_0_4 = 0;
localparam cast_sid_0_4 = 0;
localparam gather_sid_0_4 = 0;

localparam cast_out_0_5 = 0;
localparam merge_out_0_5 = 1;
localparam gather_out_0_5 = 0;
localparam merge_in_0_5 = 0;
localparam gather_in_0_5 = 0;
localparam cast_sid_0_5 = 0;
localparam gather_sid_0_5 = 0;

localparam cast_out_0_6 = 0;
localparam merge_out_0_6 = 1;
localparam gather_out_0_6 = 0;
localparam merge_in_0_6 = 0;
localparam gather_in_0_6 = 0;
localparam cast_sid_0_6 = 0;
localparam gather_sid_0_6 = 0;

localparam cast_out_0_7 = 1;
localparam merge_out_0_7 = 0;
localparam gather_out_0_7 = 0;
localparam merge_in_0_7 = 1;
localparam gather_in_0_7 = 0;
localparam cast_sid_0_7 = 19;
localparam gather_sid_0_7 = 0;

localparam cast_out_0_8 = 0;
localparam merge_out_0_8 = 1;
localparam gather_out_0_8 = 0;
localparam merge_in_0_8 = 0;
localparam gather_in_0_8 = 0;
localparam cast_sid_0_8 = 0;
localparam gather_sid_0_8 = 0;

localparam cast_out_0_9 = 0;
localparam merge_out_0_9 = 0;
localparam gather_out_0_9 = 0;
localparam merge_in_0_9 = 0;
localparam gather_in_0_9 = 0;
localparam cast_sid_0_9 = 0;
localparam gather_sid_0_9 = 0;

localparam cast_out_1_0 = 1;
localparam merge_out_1_0 = 0;
localparam gather_out_1_0 = 0;
localparam merge_in_1_0 = 0;
localparam gather_in_1_0 = 0;
localparam cast_sid_1_0 = 2;
localparam gather_sid_1_0 = 0;

localparam cast_out_1_1 = 1;
localparam merge_out_1_1 = 0;
localparam gather_out_1_1 = 0;
localparam merge_in_1_1 = 0;
localparam gather_in_1_1 = 0;
localparam cast_sid_1_1 = 8;
localparam gather_sid_1_1 = 0;

localparam cast_out_1_2 = 0;
localparam merge_out_1_2 = 0;
localparam gather_out_1_2 = 1;
localparam merge_in_1_2 = 0;
localparam gather_in_1_2 = 0;
localparam cast_sid_1_2 = 0;
localparam gather_sid_1_2 = 6;

localparam cast_out_1_3 = 0;
localparam merge_out_1_3 = 1;
localparam gather_out_1_3 = 0;
localparam merge_in_1_3 = 0;
localparam gather_in_1_3 = 0;
localparam cast_sid_1_3 = 0;
localparam gather_sid_1_3 = 0;

localparam cast_out_1_4 = 1;
localparam merge_out_1_4 = 0;
localparam gather_out_1_4 = 0;
localparam merge_in_1_4 = 1;
localparam gather_in_1_4 = 0;
localparam cast_sid_1_4 = 15;
localparam gather_sid_1_4 = 0;

localparam cast_out_1_5 = 0;
localparam merge_out_1_5 = 1;
localparam gather_out_1_5 = 0;
localparam merge_in_1_5 = 0;
localparam gather_in_1_5 = 0;
localparam cast_sid_1_5 = 0;
localparam gather_sid_1_5 = 0;

localparam cast_out_1_6 = 1;
localparam merge_out_1_6 = 0;
localparam gather_out_1_6 = 1;
localparam merge_in_1_6 = 1;
localparam gather_in_1_6 = 1;
localparam cast_sid_1_6 = 17;
localparam gather_sid_1_6 = 8;

localparam cast_out_1_7 = 0;
localparam merge_out_1_7 = 1;
localparam gather_out_1_7 = 0;
localparam merge_in_1_7 = 0;
localparam gather_in_1_7 = 0;
localparam cast_sid_1_7 = 0;
localparam gather_sid_1_7 = 0;

localparam cast_out_1_8 = 0;
localparam merge_out_1_8 = 1;
localparam gather_out_1_8 = 0;
localparam merge_in_1_8 = 0;
localparam gather_in_1_8 = 0;
localparam cast_sid_1_8 = 0;
localparam gather_sid_1_8 = 0;

localparam cast_out_1_9 = 0;
localparam merge_out_1_9 = 0;
localparam gather_out_1_9 = 0;
localparam merge_in_1_9 = 0;
localparam gather_in_1_9 = 0;
localparam cast_sid_1_9 = 0;
localparam gather_sid_1_9 = 0;

localparam cast_out_2_0 = 1;
localparam merge_out_2_0 = 0;
localparam gather_out_2_0 = 1;
localparam merge_in_2_0 = 0;
localparam gather_in_2_0 = 1;
localparam cast_sid_2_0 = 3;
localparam gather_sid_2_0 = 2;

localparam cast_out_2_1 = 1;
localparam merge_out_2_1 = 0;
localparam gather_out_2_1 = 1;
localparam merge_in_2_1 = 0;
localparam gather_in_2_1 = 1;
localparam cast_sid_2_1 = 7;
localparam gather_sid_2_1 = 3;

localparam cast_out_2_2 = 0;
localparam merge_out_2_2 = 1;
localparam gather_out_2_2 = 0;
localparam merge_in_2_2 = 0;
localparam gather_in_2_2 = 0;
localparam cast_sid_2_2 = 0;
localparam gather_sid_2_2 = 0;

localparam cast_out_2_3 = 0;
localparam merge_out_2_3 = 1;
localparam gather_out_2_3 = 0;
localparam merge_in_2_3 = 0;
localparam gather_in_2_3 = 0;
localparam cast_sid_2_3 = 0;
localparam gather_sid_2_3 = 0;

localparam cast_out_2_4 = 0;
localparam merge_out_2_4 = 0;
localparam gather_out_2_4 = 1;
localparam merge_in_2_4 = 0;
localparam gather_in_2_4 = 0;
localparam cast_sid_2_4 = 0;
localparam gather_sid_2_4 = 9;

localparam cast_out_2_5 = 1;
localparam merge_out_2_5 = 0;
localparam gather_out_2_5 = 1;
localparam merge_in_2_5 = 1;
localparam gather_in_2_5 = 1;
localparam cast_sid_2_5 = 16;
localparam gather_sid_2_5 = 7;

localparam cast_out_2_6 = 0;
localparam merge_out_2_6 = 1;
localparam gather_out_2_6 = 0;
localparam merge_in_2_6 = 0;
localparam gather_in_2_6 = 0;
localparam cast_sid_2_6 = 0;
localparam gather_sid_2_6 = 0;

localparam cast_out_2_7 = 0;
localparam merge_out_2_7 = 1;
localparam gather_out_2_7 = 0;
localparam merge_in_2_7 = 0;
localparam gather_in_2_7 = 0;
localparam cast_sid_2_7 = 0;
localparam gather_sid_2_7 = 0;

localparam cast_out_2_8 = 0;
localparam merge_out_2_8 = 1;
localparam gather_out_2_8 = 0;
localparam merge_in_2_8 = 0;
localparam gather_in_2_8 = 0;
localparam cast_sid_2_8 = 0;
localparam gather_sid_2_8 = 0;

localparam cast_out_2_9 = 0;
localparam merge_out_2_9 = 1;
localparam gather_out_2_9 = 0;
localparam merge_in_2_9 = 0;
localparam gather_in_2_9 = 0;
localparam cast_sid_2_9 = 0;
localparam gather_sid_2_9 = 0;

localparam cast_out_3_0 = 1;
localparam merge_out_3_0 = 0;
localparam gather_out_3_0 = 0;
localparam merge_in_3_0 = 0;
localparam gather_in_3_0 = 0;
localparam cast_sid_3_0 = 4;
localparam gather_sid_3_0 = 0;

localparam cast_out_3_1 = 0;
localparam merge_out_3_1 = 0;
localparam gather_out_3_1 = 1;
localparam merge_in_3_1 = 0;
localparam gather_in_3_1 = 0;
localparam cast_sid_3_1 = 0;
localparam gather_sid_3_1 = 4;

localparam cast_out_3_2 = 1;
localparam merge_out_3_2 = 0;
localparam gather_out_3_2 = 1;
localparam merge_in_3_2 = 1;
localparam gather_in_3_2 = 1;
localparam cast_sid_3_2 = 11;
localparam gather_sid_3_2 = 5;

localparam cast_out_3_3 = 1;
localparam merge_out_3_3 = 0;
localparam gather_out_3_3 = 0;
localparam merge_in_3_3 = 1;
localparam gather_in_3_3 = 1;
localparam cast_sid_3_3 = 13;
localparam gather_sid_3_3 = 0;

localparam cast_out_3_4 = 0;
localparam merge_out_3_4 = 0;
localparam gather_out_3_4 = 1;
localparam merge_in_3_4 = 0;
localparam gather_in_3_4 = 0;
localparam cast_sid_3_4 = 0;
localparam gather_sid_3_4 = 10;

localparam cast_out_3_5 = 0;
localparam merge_out_3_5 = 1;
localparam gather_out_3_5 = 0;
localparam merge_in_3_5 = 0;
localparam gather_in_3_5 = 0;
localparam cast_sid_3_5 = 0;
localparam gather_sid_3_5 = 0;

localparam cast_out_3_6 = 0;
localparam merge_out_3_6 = 1;
localparam gather_out_3_6 = 0;
localparam merge_in_3_6 = 0;
localparam gather_in_3_6 = 0;
localparam cast_sid_3_6 = 0;
localparam gather_sid_3_6 = 0;

localparam cast_out_3_7 = 0;
localparam merge_out_3_7 = 1;
localparam gather_out_3_7 = 0;
localparam merge_in_3_7 = 0;
localparam gather_in_3_7 = 0;
localparam cast_sid_3_7 = 0;
localparam gather_sid_3_7 = 0;

localparam cast_out_3_8 = 1;
localparam merge_out_3_8 = 0;
localparam gather_out_3_8 = 0;
localparam merge_in_3_8 = 1;
localparam gather_in_3_8 = 1;
localparam cast_sid_3_8 = 0;
localparam gather_sid_3_8 = 0;

localparam cast_out_3_9 = 1;
localparam merge_out_3_9 = 0;
localparam gather_out_3_9 = 0;
localparam merge_in_3_9 = 1;
localparam gather_in_3_9 = 1;
localparam cast_sid_3_9 = 0;
localparam gather_sid_3_9 = 0;

localparam cast_out_4_0 = 1;
localparam merge_out_4_0 = 0;
localparam gather_out_4_0 = 0;
localparam merge_in_4_0 = 0;
localparam gather_in_4_0 = 1;
localparam cast_sid_4_0 = 5;
localparam gather_sid_4_0 = 0;

localparam cast_out_4_1 = 1;
localparam merge_out_4_1 = 0;
localparam gather_out_4_1 = 0;
localparam merge_in_4_1 = 0;
localparam gather_in_4_1 = 0;
localparam cast_sid_4_1 = 6;
localparam gather_sid_4_1 = 0;

localparam cast_out_4_2 = 0;
localparam merge_out_4_2 = 1;
localparam gather_out_4_2 = 0;
localparam merge_in_4_2 = 0;
localparam gather_in_4_2 = 0;
localparam cast_sid_4_2 = 0;
localparam gather_sid_4_2 = 0;

localparam cast_out_4_3 = 1;
localparam merge_out_4_3 = 0;
localparam gather_out_4_3 = 0;
localparam merge_in_4_3 = 1;
localparam gather_in_4_3 = 0;
localparam cast_sid_4_3 = 12;
localparam gather_sid_4_3 = 0;

localparam cast_out_4_4 = 0;
localparam merge_out_4_4 = 1;
localparam gather_out_4_4 = 0;
localparam merge_in_4_4 = 0;
localparam gather_in_4_4 = 0;
localparam cast_sid_4_4 = 0;
localparam gather_sid_4_4 = 0;

localparam cast_out_4_5 = 0;
localparam merge_out_4_5 = 1;
localparam gather_out_4_5 = 0;
localparam merge_in_4_5 = 0;
localparam gather_in_4_5 = 0;
localparam cast_sid_4_5 = 0;
localparam gather_sid_4_5 = 0;

localparam cast_out_4_6 = 0;
localparam merge_out_4_6 = 1;
localparam gather_out_4_6 = 0;
localparam merge_in_4_6 = 0;
localparam gather_in_4_6 = 0;
localparam cast_sid_4_6 = 0;
localparam gather_sid_4_6 = 0;

localparam cast_out_4_7 = 1;
localparam merge_out_4_7 = 0;
localparam gather_out_4_7 = 0;
localparam merge_in_4_7 = 1;
localparam gather_in_4_7 = 0;
localparam cast_sid_4_7 = 18;
localparam gather_sid_4_7 = 0;

localparam cast_out_4_8 = 0;
localparam merge_out_4_8 = 1;
localparam gather_out_4_8 = 0;
localparam merge_in_4_8 = 0;
localparam gather_in_4_8 = 0;
localparam cast_sid_4_8 = 0;
localparam gather_sid_4_8 = 0;

localparam cast_out_4_9 = 0;
localparam merge_out_4_9 = 1;
localparam gather_out_4_9 = 0;
localparam merge_in_4_9 = 0;
localparam gather_in_4_9 = 0;
localparam cast_sid_4_9 = 0;
localparam gather_sid_4_9 = 0;

`endif

